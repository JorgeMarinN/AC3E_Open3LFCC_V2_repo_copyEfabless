magic
tech sky130A
timestamp 1699287058
<< checkpaint >>
rect -630 37170 25730 89430
rect -630 -630 19130 37170
<< metal2 >>
rect 3000 83060 5200 83600
rect 3000 82870 4960 83060
rect 3000 82000 5200 82870
rect 3000 42760 5740 43000
rect 5930 42760 6800 43000
rect 3000 41400 6800 42760
rect 3000 32440 6800 33800
rect 3000 32200 5740 32440
rect 5930 32200 6800 32440
rect 3000 5749 4962 6000
rect 3000 5200 5300 5749
<< metal3 >>
rect 6000 84600 23900 87600
rect 1000 67700 4000 81600
rect 20900 69700 23900 84600
rect 1000 58700 18900 67700
rect 1000 43800 4000 58700
rect 20900 41800 23900 56700
rect 6000 38800 23900 41800
rect 6000 33800 17900 38800
rect 1000 22900 4000 31800
rect 14900 24900 17900 33800
rect 1000 14900 12900 22900
rect 1000 7000 4000 14900
rect 14900 4000 17900 12900
rect 6000 1000 17900 4000
<< metal4 >>
rect 6000 84600 23900 87600
rect 1000 67700 4000 81600
rect 20900 69700 23900 84600
rect 1000 58700 18900 67700
rect 1000 43800 4000 58700
rect 20900 41800 23900 56700
rect 6000 38800 23900 41800
rect 6000 33800 17900 38800
rect 1000 22900 4000 31800
rect 14900 24900 17900 33800
rect 1000 14900 12900 22900
rect 1000 7000 4000 14900
rect 14900 4000 17900 12900
rect 6000 1000 17900 4000
<< metal5 >>
rect 6000 84600 23900 87600
rect 1000 67700 4000 81600
rect 20900 69700 23900 84600
rect 1000 58700 18900 67700
rect 1000 43800 4000 58700
rect 20900 41800 23900 56700
rect 6000 38800 23900 41800
rect 6000 33800 17900 38800
rect 1000 22900 4000 31800
rect 14900 24900 17900 33800
rect 1000 14900 12900 22900
rect 1000 7000 4000 14900
rect 14900 4000 17900 12900
rect 6000 1000 17900 4000
use nmos_waffle_14x14  nmos_waffle_14x14_0
timestamp 1699286800
transform 1 0 5925 0 1 5975
box -5925 -5975 12575 12525
use nmos_waffle_14x14  nmos_waffle_14x14_1
timestamp 1699286800
transform 0 1 5975 -1 0 31475
box -5925 -5975 12575 12525
use pmos_waffle_26x26  pmos_waffle_26x26_0
timestamp 1699286806
transform 0 1 5975 1 0 43725
box -5925 -5975 19175 19125
use pmos_waffle_26x26  pmos_waffle_26x26_1
timestamp 1699286806
transform 1 0 5925 0 -1 82825
box -5925 -5975 19175 19125
<< labels >>
rlabel metal5 6000 85600 7000 86600 7 VP
rlabel metal2 3000 82600 4000 83600 7 s1
rlabel metal5 1000 62700 2000 63700 7 fc1
rlabel metal2 3000 41800 4000 42800 7 s2
rlabel metal5 6000 36800 12500 37800 7 out
rlabel metal2 3000 32800 4000 33800 7 s3
rlabel metal5 1000 18400 2000 19400 7 fc2
rlabel metal2 3000 5500 4000 6000 7 s4
rlabel metal5 6000 2000 7000 3000 7 VN
<< end >>
