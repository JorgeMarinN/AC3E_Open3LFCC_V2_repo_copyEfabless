magic
tech sky130A
magscale 1 2
timestamp 1699299084
<< checkpaint >>
rect -3932 125824 54132 181532
rect 0 66465 54132 125824
rect -16265 -3065 193865 66465
rect -3932 -3932 193865 -3065
rect 59335 -16265 193865 -3932
<< obsactive >>
rect -12333 56652 189933 62533
rect -12333 50602 7650 56652
rect 16586 50602 61150 56652
rect 70086 50602 79650 56652
rect 88586 50602 161550 56652
rect 170486 50602 189933 56652
rect -12333 50200 189933 50602
rect -12333 13200 0 50200
rect 37000 13200 37800 50200
rect 74800 13200 75600 50200
rect -12333 867 75600 13200
rect 63267 0 75600 867
rect 125800 0 127400 50200
rect 177600 0 189933 50200
rect 63267 -12333 189933 0
<< metal1 >>
rect 2000 59000 177550 59600
rect 11150 58890 177550 58900
rect 11150 58710 11160 58890
rect 11340 58710 177550 58890
rect 11150 58700 177550 58710
rect 64650 58590 177550 58600
rect 64650 58410 64660 58590
rect 64840 58410 177550 58590
rect 64650 58400 177550 58410
rect 83150 58290 177550 58300
rect 83150 58110 83160 58290
rect 83340 58110 177550 58290
rect 83150 58100 177550 58110
rect 165050 57990 177550 58000
rect 165050 57810 165060 57990
rect 165240 57810 177550 57990
rect 165050 57800 177550 57810
rect 2000 57690 178550 57700
rect 2000 57210 10844 57690
rect 10910 57210 64344 57690
rect 64410 57210 82844 57690
rect 82910 57210 164744 57690
rect 164810 57210 178550 57690
rect 2000 57200 178550 57210
rect 2000 56500 177550 57100
<< via1 >>
rect 11160 58710 11340 58890
rect 64660 58410 64840 58590
rect 83160 58110 83340 58290
rect 165060 57810 165240 57990
rect 10844 57210 10910 57690
rect 64344 57210 64410 57690
rect 82844 57210 82910 57690
rect 164744 57210 164810 57690
rect 10844 55612 10910 56072
rect 11720 55412 11900 55992
rect 64344 55612 64410 56072
rect 65220 55412 65400 55992
rect 82844 55612 82910 56072
rect 83720 55412 83900 55992
rect 164744 55612 164810 56072
rect 165620 55412 165800 55992
<< metal2 >>
rect 5000 51790 6000 59600
rect 11150 58890 11350 58900
rect 11150 58710 11160 58890
rect 11340 58710 11350 58890
rect 10834 57690 10920 57700
rect 10834 57210 10844 57690
rect 10910 57210 10920 57690
rect 10834 56072 10920 57210
rect 11150 56332 11350 58710
rect 10834 55612 10844 56072
rect 10910 55612 10920 56072
rect 10834 55602 10920 55612
rect 11710 55992 11910 59600
rect 64650 58590 64850 58600
rect 64650 58410 64660 58590
rect 64840 58410 64850 58590
rect 11710 55412 11720 55992
rect 11900 55412 11910 55992
rect 64334 57690 64420 57700
rect 64334 57210 64344 57690
rect 64410 57210 64420 57690
rect 64334 56072 64420 57210
rect 64650 56332 64850 58410
rect 64334 55612 64344 56072
rect 64410 55612 64420 56072
rect 64334 55602 64420 55612
rect 65210 55992 65410 59600
rect 83150 58290 83350 58300
rect 83150 58110 83160 58290
rect 83340 58110 83350 58290
rect 11710 55402 11910 55412
rect 65210 55412 65220 55992
rect 65400 55412 65410 55992
rect 82834 57690 82920 57700
rect 82834 57210 82844 57690
rect 82910 57210 82920 57690
rect 82834 56072 82920 57210
rect 83150 56332 83350 58110
rect 82834 55612 82844 56072
rect 82910 55612 82920 56072
rect 82834 55602 82920 55612
rect 83710 55992 83910 59600
rect 165050 57990 165250 58000
rect 165050 57810 165060 57990
rect 165240 57810 165250 57990
rect 65210 55402 65410 55412
rect 83710 55412 83720 55992
rect 83900 55412 83910 55992
rect 164734 57690 164820 57700
rect 164734 57210 164744 57690
rect 164810 57210 164820 57690
rect 164734 56072 164820 57210
rect 165050 56332 165250 57810
rect 164734 55612 164744 56072
rect 164810 55612 164820 56072
rect 164734 55602 164820 55612
rect 165610 55992 165810 59600
rect 83710 55402 83910 55412
rect 165610 55412 165620 55992
rect 165800 55412 165810 55992
rect 165610 55402 165810 55412
rect 5000 50810 5010 51790
rect 5990 50810 6000 51790
rect 5000 50800 6000 50810
rect 172550 51790 173550 57700
rect 172550 50810 172560 51790
rect 173540 50810 173550 51790
rect 172550 50800 173550 50810
rect 11744 44572 12344 50702
rect 11744 43832 11774 44572
rect 12314 43832 12344 44572
rect 11744 43802 12344 43832
rect 65244 44572 65844 50702
rect 65244 43832 65274 44572
rect 65814 43832 65844 44572
rect 65244 43802 65844 43832
rect 83744 44572 84344 50702
rect 83744 43832 83774 44572
rect 84314 43832 84344 44572
rect 83744 43802 84344 43832
rect 165644 44572 166244 50702
rect 165644 43832 165674 44572
rect 166214 43832 166244 44572
rect 165644 43802 166244 43832
<< via2 >>
rect 5010 50810 5990 51790
rect 172560 50810 173540 51790
rect 11774 43832 12314 44572
rect 65274 43832 65814 44572
rect 83774 43832 84314 44572
rect 165674 43832 166214 44572
<< metal3 >>
rect 5000 51790 6000 51800
rect 5000 50810 5010 51790
rect 5990 50810 6000 51790
rect 5000 37800 6000 50810
rect 172550 51790 173550 51800
rect 172550 50810 172560 51790
rect 173540 50810 173550 51790
rect 11744 44572 12344 50702
rect 11744 43832 11774 44572
rect 12314 43832 12344 44572
rect 11744 43802 12344 43832
rect 65244 44572 65844 50702
rect 65244 43832 65274 44572
rect 65814 43832 65844 44572
rect 65244 43802 65844 43832
rect 83744 44572 84344 50702
rect 83744 43832 83774 44572
rect 84314 43832 84344 44572
rect 83744 43802 84344 43832
rect 165644 44572 166244 50702
rect 165644 43832 165674 44572
rect 166214 43832 166244 44572
rect 165644 43802 166244 43832
rect 172550 37800 173550 50810
<< via3 >>
rect 11774 43832 12314 44572
rect 65274 43832 65814 44572
rect 83774 43832 84314 44572
rect 165674 43832 166214 44572
<< metal4 >>
rect 11744 44572 12344 50702
rect 11744 43832 11774 44572
rect 12314 43832 12344 44572
rect 11744 43802 12344 43832
rect 65244 44572 65844 50702
rect 65244 43832 65274 44572
rect 65814 43832 65844 44572
rect 65244 43802 65844 43832
rect 83744 44572 84344 50702
rect 83744 43832 83774 44572
rect 84314 43832 84344 44572
rect 83744 43802 84344 43832
rect 165644 44572 166244 50702
rect 165644 43832 165674 44572
rect 166214 43832 166244 44572
rect 165644 43802 166244 43832
<< via4 >>
rect 11774 43832 12314 44572
rect 65274 43832 65814 44572
rect 83774 43832 84314 44572
rect 165674 43832 166214 44572
<< metal5 >>
rect 11744 44572 12344 50702
rect 11744 43832 11774 44572
rect 12314 43832 12344 44572
rect 11744 43802 12344 43832
rect 65244 44572 65844 50702
rect 65244 43832 65274 44572
rect 65814 43832 65844 44572
rect 65244 43802 65844 43832
rect 83744 44572 84344 50702
rect 83744 43832 83774 44572
rect 84314 43832 84344 44572
rect 83744 43802 84344 43832
rect 165644 44572 166244 50702
rect 165644 43832 165674 44572
rect 166214 43832 166244 44572
rect 165644 43802 166244 43832
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 161550 -1 0 56652
box 0 0 6050 8936
use level_shifter  level_shifter_1
timestamp 1666543010
transform 0 1 79650 -1 0 56652
box 0 0 6050 8936
use level_shifter  level_shifter_2
timestamp 1666543010
transform 0 1 61150 -1 0 56652
box 0 0 6050 8936
use level_shifter  level_shifter_3
timestamp 1666543010
transform 0 1 7650 -1 0 56652
box 0 0 6050 8936
use power_stage_2  power_stage_2_0
timestamp 1699287058
transform 0 1 0 -1 0 50200
box 0 0 50200 177600
<< labels >>
rlabel metal1 164350 56500 177550 57100 3 VLS
rlabel metal1 165350 57200 178550 57700 7 VDD
rlabel metal1 177350 57800 177550 58000 7 D1
rlabel metal1 177350 58100 177550 58300 7 D2
rlabel metal1 177350 58400 177550 58600 7 D3
rlabel metal1 177350 58700 177550 58900 7 D4
<< end >>
