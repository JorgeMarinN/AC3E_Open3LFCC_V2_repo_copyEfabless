magic
tech sky130A
magscale 1 2
timestamp 1700268818
<< nwell >>
rect 221 954 3483 2502
rect -395 88 3483 954
<< mvnmos >>
rect -129 -754 -29 -154
rect 29 -754 129 -154
rect 459 -954 559 -154
rect 617 -954 717 -154
rect 775 -954 875 -154
rect 933 -954 1033 -154
rect 1091 -954 1191 -154
rect 1249 -954 1349 -154
rect 1407 -954 1507 -154
rect 1565 -954 1665 -154
rect 1723 -954 1823 -154
rect 1881 -954 1981 -154
rect 2039 -954 2139 -154
rect 2197 -954 2297 -154
rect 2355 -954 2455 -154
rect 2513 -954 2613 -154
rect 2671 -954 2771 -154
rect 2829 -954 2929 -154
rect 2987 -954 3087 -154
rect 3145 -954 3245 -154
<< mvpmos >>
rect -137 154 -37 354
rect 37 154 137 754
rect 459 154 559 2322
rect 617 154 717 2322
rect 775 154 875 2322
rect 933 154 1033 2322
rect 1091 154 1191 2322
rect 1249 154 1349 2322
rect 1407 154 1507 2322
rect 1565 154 1665 2322
rect 1723 154 1823 2322
rect 1881 154 1981 2322
rect 2039 154 2139 2322
rect 2197 154 2297 2322
rect 2355 154 2455 2322
rect 2513 154 2613 2322
rect 2671 154 2771 2322
rect 2829 154 2929 2322
rect 2987 154 3087 2322
rect 3145 154 3245 2322
<< mvndiff >>
rect -187 -166 -129 -154
rect -187 -742 -175 -166
rect -141 -742 -129 -166
rect -187 -754 -129 -742
rect -29 -166 29 -154
rect -29 -742 -17 -166
rect 17 -742 29 -166
rect -29 -754 29 -742
rect 129 -166 187 -154
rect 129 -742 141 -166
rect 175 -742 187 -166
rect 129 -754 187 -742
rect 401 -166 459 -154
rect 401 -942 413 -166
rect 447 -942 459 -166
rect 401 -954 459 -942
rect 559 -166 617 -154
rect 559 -942 571 -166
rect 605 -942 617 -166
rect 559 -954 617 -942
rect 717 -166 775 -154
rect 717 -942 729 -166
rect 763 -942 775 -166
rect 717 -954 775 -942
rect 875 -166 933 -154
rect 875 -942 887 -166
rect 921 -942 933 -166
rect 875 -954 933 -942
rect 1033 -166 1091 -154
rect 1033 -942 1045 -166
rect 1079 -942 1091 -166
rect 1033 -954 1091 -942
rect 1191 -166 1249 -154
rect 1191 -942 1203 -166
rect 1237 -942 1249 -166
rect 1191 -954 1249 -942
rect 1349 -166 1407 -154
rect 1349 -942 1361 -166
rect 1395 -942 1407 -166
rect 1349 -954 1407 -942
rect 1507 -166 1565 -154
rect 1507 -942 1519 -166
rect 1553 -942 1565 -166
rect 1507 -954 1565 -942
rect 1665 -166 1723 -154
rect 1665 -942 1677 -166
rect 1711 -942 1723 -166
rect 1665 -954 1723 -942
rect 1823 -166 1881 -154
rect 1823 -942 1835 -166
rect 1869 -942 1881 -166
rect 1823 -954 1881 -942
rect 1981 -166 2039 -154
rect 1981 -942 1993 -166
rect 2027 -942 2039 -166
rect 1981 -954 2039 -942
rect 2139 -166 2197 -154
rect 2139 -942 2151 -166
rect 2185 -942 2197 -166
rect 2139 -954 2197 -942
rect 2297 -166 2355 -154
rect 2297 -942 2309 -166
rect 2343 -942 2355 -166
rect 2297 -954 2355 -942
rect 2455 -166 2513 -154
rect 2455 -942 2467 -166
rect 2501 -942 2513 -166
rect 2455 -954 2513 -942
rect 2613 -166 2671 -154
rect 2613 -942 2625 -166
rect 2659 -942 2671 -166
rect 2613 -954 2671 -942
rect 2771 -166 2829 -154
rect 2771 -942 2783 -166
rect 2817 -942 2829 -166
rect 2771 -954 2829 -942
rect 2929 -166 2987 -154
rect 2929 -942 2941 -166
rect 2975 -942 2987 -166
rect 2929 -954 2987 -942
rect 3087 -166 3145 -154
rect 3087 -942 3099 -166
rect 3133 -942 3145 -166
rect 3087 -954 3145 -942
rect 3245 -166 3303 -154
rect 3245 -942 3257 -166
rect 3291 -942 3303 -166
rect 3245 -954 3303 -942
<< mvpdiff >>
rect -21 742 37 754
rect -21 354 -9 742
rect -195 342 -137 354
rect -195 166 -183 342
rect -149 166 -137 342
rect -195 154 -137 166
rect -37 342 -9 354
rect -37 166 -25 342
rect 25 166 37 742
rect -37 154 37 166
rect 137 742 195 754
rect 137 166 149 742
rect 183 166 195 742
rect 137 154 195 166
rect 401 2310 459 2322
rect 401 166 413 2310
rect 447 166 459 2310
rect 401 154 459 166
rect 559 2310 617 2322
rect 559 166 571 2310
rect 605 166 617 2310
rect 559 154 617 166
rect 717 2310 775 2322
rect 717 166 729 2310
rect 763 166 775 2310
rect 717 154 775 166
rect 875 2310 933 2322
rect 875 166 887 2310
rect 921 166 933 2310
rect 875 154 933 166
rect 1033 2310 1091 2322
rect 1033 166 1045 2310
rect 1079 166 1091 2310
rect 1033 154 1091 166
rect 1191 2310 1249 2322
rect 1191 166 1203 2310
rect 1237 166 1249 2310
rect 1191 154 1249 166
rect 1349 2310 1407 2322
rect 1349 166 1361 2310
rect 1395 166 1407 2310
rect 1349 154 1407 166
rect 1507 2310 1565 2322
rect 1507 166 1519 2310
rect 1553 166 1565 2310
rect 1507 154 1565 166
rect 1665 2310 1723 2322
rect 1665 166 1677 2310
rect 1711 166 1723 2310
rect 1665 154 1723 166
rect 1823 2310 1881 2322
rect 1823 166 1835 2310
rect 1869 166 1881 2310
rect 1823 154 1881 166
rect 1981 2310 2039 2322
rect 1981 166 1993 2310
rect 2027 166 2039 2310
rect 1981 154 2039 166
rect 2139 2310 2197 2322
rect 2139 166 2151 2310
rect 2185 166 2197 2310
rect 2139 154 2197 166
rect 2297 2310 2355 2322
rect 2297 166 2309 2310
rect 2343 166 2355 2310
rect 2297 154 2355 166
rect 2455 2310 2513 2322
rect 2455 166 2467 2310
rect 2501 166 2513 2310
rect 2455 154 2513 166
rect 2613 2310 2671 2322
rect 2613 166 2625 2310
rect 2659 166 2671 2310
rect 2613 154 2671 166
rect 2771 2310 2829 2322
rect 2771 166 2783 2310
rect 2817 166 2829 2310
rect 2771 154 2829 166
rect 2929 2310 2987 2322
rect 2929 166 2941 2310
rect 2975 166 2987 2310
rect 2929 154 2987 166
rect 3087 2310 3145 2322
rect 3087 166 3099 2310
rect 3133 166 3145 2310
rect 3087 154 3145 166
rect 3245 2310 3303 2322
rect 3245 166 3257 2310
rect 3291 166 3303 2310
rect 3245 154 3303 166
<< mvndiffc >>
rect -175 -742 -141 -166
rect -17 -742 17 -166
rect 141 -742 175 -166
rect 413 -942 447 -166
rect 571 -942 605 -166
rect 729 -942 763 -166
rect 887 -942 921 -166
rect 1045 -942 1079 -166
rect 1203 -942 1237 -166
rect 1361 -942 1395 -166
rect 1519 -942 1553 -166
rect 1677 -942 1711 -166
rect 1835 -942 1869 -166
rect 1993 -942 2027 -166
rect 2151 -942 2185 -166
rect 2309 -942 2343 -166
rect 2467 -942 2501 -166
rect 2625 -942 2659 -166
rect 2783 -942 2817 -166
rect 2941 -942 2975 -166
rect 3099 -942 3133 -166
rect 3257 -942 3291 -166
<< mvpdiffc >>
rect -183 166 -149 342
rect -9 342 25 742
rect -25 166 25 342
rect 149 166 183 742
rect 413 166 447 2310
rect 571 166 605 2310
rect 729 166 763 2310
rect 887 166 921 2310
rect 1045 166 1079 2310
rect 1203 166 1237 2310
rect 1361 166 1395 2310
rect 1519 166 1553 2310
rect 1677 166 1711 2310
rect 1835 166 1869 2310
rect 1993 166 2027 2310
rect 2151 166 2185 2310
rect 2309 166 2343 2310
rect 2467 166 2501 2310
rect 2625 166 2659 2310
rect 2783 166 2817 2310
rect 2941 166 2975 2310
rect 3099 166 3133 2310
rect 3257 166 3291 2310
<< mvpsubdiff >>
rect -301 -184 -261 -154
rect -301 -754 -261 -724
rect 287 -184 327 -154
rect -301 -982 -267 -942
rect 157 -982 187 -942
rect 287 -954 327 -924
rect 3377 -184 3417 -154
rect 3377 -954 3417 -924
rect 287 -1068 321 -1028
rect 3383 -1068 3417 -1028
<< mvnsubdiff >>
rect 307 2376 341 2416
rect 3363 2376 3397 2416
rect 307 2292 347 2322
rect -309 808 -275 848
rect 165 808 195 848
rect -289 724 -249 754
rect -289 154 -249 184
rect 307 154 347 184
rect 3357 2292 3397 2322
rect 3357 154 3397 184
<< mvpsubdiffcont >>
rect -301 -724 -261 -184
rect 287 -924 327 -184
rect -267 -982 157 -942
rect 3377 -924 3417 -184
rect 321 -1068 3383 -1028
<< mvnsubdiffcont >>
rect 341 2376 3363 2416
rect -275 808 165 848
rect -289 184 -249 724
rect 307 184 347 2292
rect 3357 184 3397 2292
<< poly >>
rect 459 2322 559 2348
rect 617 2322 717 2348
rect 775 2322 875 2348
rect 933 2322 1033 2348
rect 1091 2322 1191 2348
rect 1249 2322 1349 2348
rect 1407 2322 1507 2348
rect 1565 2322 1665 2348
rect 1723 2322 1823 2348
rect 1881 2322 1981 2348
rect 2039 2322 2139 2348
rect 2197 2322 2297 2348
rect 2355 2322 2455 2348
rect 2513 2322 2613 2348
rect 2671 2322 2771 2348
rect 2829 2322 2929 2348
rect 2987 2322 3087 2348
rect 3145 2322 3245 2348
rect 37 754 137 780
rect -137 354 -37 380
rect -137 96 -37 154
rect -137 36 -117 96
rect -57 36 -37 96
rect -137 16 -37 36
rect 37 96 137 154
rect 37 36 57 96
rect 117 36 137 96
rect 37 16 137 36
rect 459 -14 559 154
rect 435 -34 559 -14
rect 435 -94 455 -34
rect 515 -94 559 -34
rect 435 -114 559 -94
rect -129 -154 -29 -128
rect 29 -154 129 -128
rect 459 -154 559 -114
rect 617 -14 717 154
rect 775 -14 875 154
rect 617 -34 875 -14
rect 617 -94 661 -34
rect 831 -94 875 -34
rect 617 -114 875 -94
rect 617 -154 717 -114
rect 775 -154 875 -114
rect 933 -14 1033 154
rect 1091 -14 1191 154
rect 933 -34 1191 -14
rect 933 -94 977 -34
rect 1147 -94 1191 -34
rect 933 -114 1191 -94
rect 933 -154 1033 -114
rect 1091 -154 1191 -114
rect 1249 -14 1349 154
rect 1407 -14 1507 154
rect 1249 -34 1507 -14
rect 1249 -94 1293 -34
rect 1463 -94 1507 -34
rect 1249 -114 1507 -94
rect 1249 -154 1349 -114
rect 1407 -154 1507 -114
rect 1565 -14 1665 154
rect 1723 -14 1823 154
rect 1565 -34 1823 -14
rect 1565 -94 1609 -34
rect 1779 -94 1823 -34
rect 1565 -114 1823 -94
rect 1565 -154 1665 -114
rect 1723 -154 1823 -114
rect 1881 -14 1981 154
rect 2039 -14 2139 154
rect 1881 -34 2139 -14
rect 1881 -94 1925 -34
rect 2095 -94 2139 -34
rect 1881 -114 2139 -94
rect 1881 -154 1981 -114
rect 2039 -154 2139 -114
rect 2197 -14 2297 154
rect 2355 -14 2455 154
rect 2197 -34 2455 -14
rect 2197 -94 2241 -34
rect 2411 -94 2455 -34
rect 2197 -114 2455 -94
rect 2197 -154 2297 -114
rect 2355 -154 2455 -114
rect 2513 -14 2613 154
rect 2671 -14 2771 154
rect 2513 -34 2771 -14
rect 2513 -94 2557 -34
rect 2727 -94 2771 -34
rect 2513 -114 2771 -94
rect 2513 -154 2613 -114
rect 2671 -154 2771 -114
rect 2829 -14 2929 154
rect 2987 -14 3087 154
rect 2829 -34 3087 -14
rect 2829 -94 2873 -34
rect 3043 -94 3087 -34
rect 2829 -114 3087 -94
rect 2829 -154 2929 -114
rect 2987 -154 3087 -114
rect 3145 -14 3245 154
rect 3145 -34 3269 -14
rect 3145 -94 3189 -34
rect 3249 -94 3269 -34
rect 3145 -114 3269 -94
rect 3145 -154 3245 -114
rect -129 -812 -29 -754
rect -129 -872 -109 -812
rect -49 -872 -29 -812
rect -129 -892 -29 -872
rect 29 -812 129 -754
rect 29 -872 49 -812
rect 109 -872 129 -812
rect 29 -892 129 -872
rect 459 -980 559 -954
rect 617 -980 717 -954
rect 775 -980 875 -954
rect 933 -980 1033 -954
rect 1091 -980 1191 -954
rect 1249 -980 1349 -954
rect 1407 -980 1507 -954
rect 1565 -980 1665 -954
rect 1723 -980 1823 -954
rect 1881 -980 1981 -954
rect 2039 -980 2139 -954
rect 2197 -980 2297 -954
rect 2355 -980 2455 -954
rect 2513 -980 2613 -954
rect 2671 -980 2771 -954
rect 2829 -980 2929 -954
rect 2987 -980 3087 -954
rect 3145 -980 3245 -954
<< polycont >>
rect -117 36 -57 96
rect 57 36 117 96
rect 455 -94 515 -34
rect 661 -94 831 -34
rect 977 -94 1147 -34
rect 1293 -94 1463 -34
rect 1609 -94 1779 -34
rect 1925 -94 2095 -34
rect 2241 -94 2411 -34
rect 2557 -94 2727 -34
rect 2873 -94 3043 -34
rect 3189 -94 3249 -34
rect -109 -872 -49 -812
rect 49 -872 109 -812
<< locali >>
rect 307 2376 341 2416
rect 3363 2376 3397 2416
rect 307 2292 347 2322
rect -309 808 -275 848
rect 165 808 195 848
rect -289 724 -249 754
rect -9 742 25 758
rect -289 154 -249 184
rect -183 342 -149 358
rect -183 150 -149 166
rect -25 342 -9 358
rect -25 150 25 166
rect 149 742 183 758
rect 149 150 183 166
rect 307 154 347 184
rect 413 2310 447 2326
rect 413 150 447 166
rect 571 2310 605 2326
rect 571 150 605 166
rect 729 2310 763 2326
rect 729 150 763 166
rect 887 2310 921 2326
rect 887 150 921 166
rect 1045 2310 1079 2326
rect 1045 150 1079 166
rect 1203 2310 1237 2326
rect 1203 150 1237 166
rect 1361 2310 1395 2326
rect 1361 150 1395 166
rect 1519 2310 1553 2326
rect 1519 150 1553 166
rect 1677 2310 1711 2326
rect 1677 150 1711 166
rect 1835 2310 1869 2326
rect 1835 150 1869 166
rect 1993 2310 2027 2326
rect 1993 150 2027 166
rect 2151 2310 2185 2326
rect 2151 150 2185 166
rect 2309 2310 2343 2326
rect 2309 150 2343 166
rect 2467 2310 2501 2326
rect 2467 150 2501 166
rect 2625 2310 2659 2326
rect 2625 150 2659 166
rect 2783 2310 2817 2326
rect 2783 150 2817 166
rect 2941 2310 2975 2326
rect 2941 150 2975 166
rect 3099 2310 3133 2326
rect 3099 150 3133 166
rect 3257 2310 3291 2326
rect 3257 150 3291 166
rect 3357 2292 3397 2322
rect 3357 154 3397 184
rect -137 96 -37 116
rect -137 36 -117 96
rect -57 36 -37 96
rect -137 -16 -37 36
rect 7 96 137 116
rect 7 36 27 96
rect 117 36 137 96
rect 7 16 137 36
rect -137 -36 -7 -16
rect -137 -96 -87 -36
rect -27 -96 -7 -36
rect -137 -116 -7 -96
rect 435 -34 535 -14
rect 435 -94 455 -34
rect 515 -94 535 -34
rect 435 -114 535 -94
rect 641 -34 851 -14
rect 641 -94 661 -34
rect 831 -94 851 -34
rect 641 -114 851 -94
rect 957 -34 1167 -14
rect 957 -94 977 -34
rect 1147 -94 1167 -34
rect 957 -114 1167 -94
rect 1273 -34 1483 -14
rect 1273 -94 1293 -34
rect 1463 -94 1483 -34
rect 1273 -114 1483 -94
rect 1589 -34 1799 -14
rect 1589 -94 1609 -34
rect 1779 -94 1799 -34
rect 1589 -114 1799 -94
rect 1905 -34 2115 -14
rect 1905 -94 1925 -34
rect 2095 -94 2115 -34
rect 1905 -114 2115 -94
rect 2221 -34 2431 -14
rect 2221 -94 2241 -34
rect 2411 -94 2431 -34
rect 2221 -114 2431 -94
rect 2537 -34 2747 -14
rect 2537 -94 2557 -34
rect 2727 -94 2747 -34
rect 2537 -114 2747 -94
rect 2853 -34 3063 -14
rect 2853 -94 2873 -34
rect 3043 -94 3063 -34
rect 2853 -114 3063 -94
rect 3169 -34 3269 -14
rect 3169 -94 3189 -34
rect 3249 -94 3269 -34
rect 3169 -114 3269 -94
rect -301 -184 -261 -154
rect -301 -754 -261 -724
rect -175 -166 -141 -150
rect -175 -758 -141 -742
rect -17 -166 17 -150
rect -17 -758 17 -742
rect 141 -166 175 -150
rect 141 -758 175 -742
rect 287 -184 327 -154
rect -151 -812 -29 -792
rect -151 -872 -131 -812
rect -49 -872 -29 -812
rect -151 -892 -29 -872
rect 29 -812 151 -792
rect 29 -872 49 -812
rect 131 -872 151 -812
rect 29 -892 151 -872
rect -301 -982 -267 -942
rect 157 -982 187 -942
rect 287 -954 327 -924
rect 413 -166 447 -150
rect 413 -958 447 -942
rect 571 -166 605 -150
rect 571 -958 605 -942
rect 729 -166 763 -150
rect 729 -958 763 -942
rect 887 -166 921 -150
rect 887 -958 921 -942
rect 1045 -166 1079 -150
rect 1045 -958 1079 -942
rect 1203 -166 1237 -150
rect 1203 -958 1237 -942
rect 1361 -166 1395 -150
rect 1361 -958 1395 -942
rect 1519 -166 1553 -150
rect 1519 -958 1553 -942
rect 1677 -166 1711 -150
rect 1677 -958 1711 -942
rect 1835 -166 1869 -150
rect 1835 -958 1869 -942
rect 1993 -166 2027 -150
rect 1993 -958 2027 -942
rect 2151 -166 2185 -150
rect 2151 -958 2185 -942
rect 2309 -166 2343 -150
rect 2309 -958 2343 -942
rect 2467 -166 2501 -150
rect 2467 -958 2501 -942
rect 2625 -166 2659 -150
rect 2625 -958 2659 -942
rect 2783 -166 2817 -150
rect 2783 -958 2817 -942
rect 2941 -166 2975 -150
rect 2941 -958 2975 -942
rect 3099 -166 3133 -150
rect 3099 -958 3133 -942
rect 3257 -166 3291 -150
rect 3257 -958 3291 -942
rect 3377 -184 3417 -154
rect 3377 -954 3417 -924
rect 287 -1068 321 -1028
rect 3383 -1068 3417 -1028
<< viali >>
rect 341 2376 3363 2416
rect -275 808 165 848
rect -289 184 -249 724
rect -183 166 -149 342
rect -9 342 25 742
rect -25 166 25 342
rect 149 166 183 742
rect 307 184 347 2292
rect 413 166 447 2310
rect 571 166 605 2310
rect 729 166 763 2310
rect 887 166 921 2310
rect 1045 166 1079 2310
rect 1203 166 1237 2310
rect 1361 166 1395 2310
rect 1519 166 1553 2310
rect 1677 166 1711 2310
rect 1835 166 1869 2310
rect 1993 166 2027 2310
rect 2151 166 2185 2310
rect 2309 166 2343 2310
rect 2467 166 2501 2310
rect 2625 166 2659 2310
rect 2783 166 2817 2310
rect 2941 166 2975 2310
rect 3099 166 3133 2310
rect 3257 166 3291 2310
rect 3357 184 3397 2292
rect 27 36 57 96
rect 57 36 87 96
rect -87 -96 -27 -36
rect 455 -94 515 -34
rect 661 -94 831 -34
rect 977 -94 1147 -34
rect 1293 -94 1463 -34
rect 1609 -94 1779 -34
rect 1925 -94 2095 -34
rect 2241 -94 2411 -34
rect 2557 -94 2727 -34
rect 2873 -94 3043 -34
rect 3189 -94 3249 -34
rect -301 -724 -261 -184
rect -175 -742 -141 -166
rect -17 -742 17 -166
rect 141 -742 175 -166
rect -131 -872 -109 -812
rect -109 -872 -71 -812
rect 71 -872 109 -812
rect 109 -872 131 -812
rect 287 -924 327 -184
rect -267 -982 157 -942
rect 413 -942 447 -166
rect 571 -942 605 -166
rect 729 -942 763 -166
rect 887 -942 921 -166
rect 1045 -942 1079 -166
rect 1203 -942 1237 -166
rect 1361 -942 1395 -166
rect 1519 -942 1553 -166
rect 1677 -942 1711 -166
rect 1835 -942 1869 -166
rect 1993 -942 2027 -166
rect 2151 -942 2185 -166
rect 2309 -942 2343 -166
rect 2467 -942 2501 -166
rect 2625 -942 2659 -166
rect 2783 -942 2817 -166
rect 2941 -942 2975 -166
rect 3099 -942 3133 -166
rect 3257 -942 3291 -166
rect 3377 -924 3417 -184
rect 321 -1068 3383 -1028
<< metal1 >>
rect 287 2416 3417 2436
rect 287 2376 341 2416
rect 3363 2376 3417 2416
rect 287 2356 3417 2376
rect 287 2310 453 2356
rect 287 2292 413 2310
rect 287 988 307 2292
rect -309 848 307 988
rect -309 808 -275 848
rect 165 808 307 848
rect -309 788 307 808
rect -309 724 -229 788
rect -309 184 -289 724
rect -249 184 -229 724
rect -15 742 31 788
rect -15 354 -9 742
rect -309 154 -229 184
rect -189 342 -143 354
rect -189 166 -183 342
rect -149 166 -143 342
rect -189 116 -143 166
rect -31 342 -9 354
rect -31 166 -25 342
rect 25 166 31 742
rect -31 154 31 166
rect 143 742 189 754
rect 143 166 149 742
rect 183 166 189 742
rect -189 96 107 116
rect -189 36 27 96
rect 87 36 107 96
rect -189 16 107 36
rect -321 -184 -241 -154
rect -321 -724 -301 -184
rect -261 -724 -241 -184
rect -321 -922 -241 -724
rect -181 -166 -135 16
rect 143 -16 189 166
rect 287 184 307 788
rect 347 184 413 2292
rect 287 166 413 184
rect 447 166 453 2310
rect 287 154 453 166
rect 565 2310 611 2322
rect 565 166 571 2310
rect 605 166 611 2310
rect 565 114 611 166
rect 723 2310 769 2356
rect 723 166 729 2310
rect 763 166 769 2310
rect 723 154 769 166
rect 881 2310 927 2322
rect 881 166 887 2310
rect 921 166 927 2310
rect 881 114 927 166
rect 1039 2310 1085 2356
rect 1039 166 1045 2310
rect 1079 166 1085 2310
rect 1039 154 1085 166
rect 1197 2310 1243 2322
rect 1197 166 1203 2310
rect 1237 166 1243 2310
rect 1197 114 1243 166
rect 1355 2310 1401 2356
rect 1355 166 1361 2310
rect 1395 166 1401 2310
rect 1355 154 1401 166
rect 1513 2310 1559 2322
rect 1513 166 1519 2310
rect 1553 166 1559 2310
rect 1513 114 1559 166
rect 1671 2310 1717 2356
rect 1671 166 1677 2310
rect 1711 166 1717 2310
rect 1671 154 1717 166
rect 1829 2310 1875 2322
rect 1829 166 1835 2310
rect 1869 166 1875 2310
rect 1829 114 1875 166
rect 1987 2310 2033 2356
rect 1987 166 1993 2310
rect 2027 166 2033 2310
rect 1987 154 2033 166
rect 2145 2310 2191 2322
rect 2145 166 2151 2310
rect 2185 166 2191 2310
rect 2145 114 2191 166
rect 2303 2310 2349 2356
rect 2303 166 2309 2310
rect 2343 166 2349 2310
rect 2303 154 2349 166
rect 2461 2310 2507 2322
rect 2461 166 2467 2310
rect 2501 166 2507 2310
rect 2461 114 2507 166
rect 2619 2310 2665 2356
rect 2619 166 2625 2310
rect 2659 166 2665 2310
rect 2619 154 2665 166
rect 2777 2310 2823 2322
rect 2777 166 2783 2310
rect 2817 166 2823 2310
rect 2777 114 2823 166
rect 2935 2310 2981 2356
rect 2935 166 2941 2310
rect 2975 166 2981 2310
rect 2935 154 2981 166
rect 3093 2310 3139 2322
rect 3093 166 3099 2310
rect 3133 166 3139 2310
rect 3093 114 3139 166
rect 3251 2310 3417 2356
rect 3251 166 3257 2310
rect 3291 2292 3417 2310
rect 3291 184 3357 2292
rect 3397 184 3417 2292
rect 3291 166 3417 184
rect 3251 154 3417 166
rect 565 94 3139 114
rect 565 34 585 94
rect 3119 34 3139 94
rect 565 14 3139 34
rect -107 -36 189 -16
rect -107 -96 -87 -36
rect -27 -96 127 -36
rect 187 -96 189 -36
rect -107 -116 189 -96
rect 435 -34 535 -14
rect 435 -94 455 -34
rect 515 -94 535 -34
rect 435 -114 535 -94
rect -181 -742 -175 -166
rect -141 -742 -135 -166
rect -181 -754 -135 -742
rect -23 -166 23 -154
rect -23 -742 -17 -166
rect 17 -742 23 -166
rect -151 -812 -51 -792
rect -151 -872 -131 -812
rect -71 -872 -51 -812
rect -151 -892 -51 -872
rect -23 -922 23 -742
rect 135 -166 181 -116
rect 135 -742 141 -166
rect 175 -742 181 -166
rect 135 -754 181 -742
rect 267 -166 453 -154
rect 267 -184 413 -166
rect 51 -812 151 -792
rect 51 -872 71 -812
rect 131 -872 151 -812
rect 51 -892 151 -872
rect 267 -922 287 -184
rect -321 -924 287 -922
rect 327 -924 413 -184
rect -321 -942 413 -924
rect 447 -942 453 -166
rect -321 -982 -267 -942
rect 157 -982 453 -942
rect 565 -166 611 14
rect 641 -34 851 -14
rect 641 -94 661 -34
rect 831 -94 851 -34
rect 641 -114 851 -94
rect 565 -942 571 -166
rect 605 -942 611 -166
rect 565 -954 611 -942
rect 723 -166 769 -154
rect 723 -942 729 -166
rect 763 -942 769 -166
rect -321 -1002 453 -982
rect 267 -1008 453 -1002
rect 723 -1008 769 -942
rect 881 -166 927 14
rect 957 -34 1167 -14
rect 957 -94 977 -34
rect 1147 -94 1167 -34
rect 957 -114 1167 -94
rect 881 -942 887 -166
rect 921 -942 927 -166
rect 881 -954 927 -942
rect 1039 -166 1085 -154
rect 1039 -942 1045 -166
rect 1079 -942 1085 -166
rect 1039 -1008 1085 -942
rect 1197 -166 1243 14
rect 1273 -34 1483 -14
rect 1273 -94 1293 -34
rect 1463 -94 1483 -34
rect 1273 -114 1483 -94
rect 1197 -942 1203 -166
rect 1237 -942 1243 -166
rect 1197 -954 1243 -942
rect 1355 -166 1401 -154
rect 1355 -942 1361 -166
rect 1395 -942 1401 -166
rect 1355 -1008 1401 -942
rect 1513 -166 1559 14
rect 1589 -34 1799 -14
rect 1589 -94 1609 -34
rect 1779 -94 1799 -34
rect 1589 -114 1799 -94
rect 1513 -942 1519 -166
rect 1553 -942 1559 -166
rect 1513 -954 1559 -942
rect 1671 -166 1717 -154
rect 1671 -942 1677 -166
rect 1711 -942 1717 -166
rect 1671 -1008 1717 -942
rect 1829 -166 1875 14
rect 1905 -34 2115 -14
rect 1905 -94 1925 -34
rect 2095 -94 2115 -34
rect 1905 -114 2115 -94
rect 1829 -942 1835 -166
rect 1869 -942 1875 -166
rect 1829 -954 1875 -942
rect 1987 -166 2033 -154
rect 1987 -942 1993 -166
rect 2027 -942 2033 -166
rect 1987 -1008 2033 -942
rect 2145 -166 2191 14
rect 2221 -34 2431 -14
rect 2221 -94 2241 -34
rect 2411 -94 2431 -34
rect 2221 -114 2431 -94
rect 2145 -942 2151 -166
rect 2185 -942 2191 -166
rect 2145 -954 2191 -942
rect 2303 -166 2349 -154
rect 2303 -942 2309 -166
rect 2343 -942 2349 -166
rect 2303 -1008 2349 -942
rect 2461 -166 2507 14
rect 2537 -34 2747 -14
rect 2537 -94 2557 -34
rect 2727 -94 2747 -34
rect 2537 -114 2747 -94
rect 2461 -942 2467 -166
rect 2501 -942 2507 -166
rect 2461 -954 2507 -942
rect 2619 -166 2665 -154
rect 2619 -942 2625 -166
rect 2659 -942 2665 -166
rect 2619 -1008 2665 -942
rect 2777 -166 2823 14
rect 2853 -34 3063 -14
rect 2853 -94 2873 -34
rect 3043 -94 3063 -34
rect 2853 -114 3063 -94
rect 2777 -942 2783 -166
rect 2817 -942 2823 -166
rect 2777 -954 2823 -942
rect 2935 -166 2981 -154
rect 2935 -942 2941 -166
rect 2975 -942 2981 -166
rect 2935 -1008 2981 -942
rect 3093 -166 3139 14
rect 3169 -34 3269 -14
rect 3169 -94 3189 -34
rect 3249 -94 3269 -34
rect 3169 -114 3269 -94
rect 3093 -942 3099 -166
rect 3133 -942 3139 -166
rect 3093 -954 3139 -942
rect 3251 -166 3437 -154
rect 3251 -942 3257 -166
rect 3291 -184 3437 -166
rect 3291 -924 3377 -184
rect 3417 -924 3437 -184
rect 3291 -942 3437 -924
rect 3251 -1008 3437 -942
rect 267 -1028 3437 -1008
rect 267 -1068 321 -1028
rect 3383 -1068 3437 -1028
rect 267 -1088 3437 -1068
<< via1 >>
rect 585 34 3119 94
rect 127 -96 187 -36
rect 455 -94 515 -34
rect -131 -872 -71 -812
rect 71 -872 131 -812
rect 661 -94 831 -34
rect 977 -94 1147 -34
rect 1293 -94 1463 -34
rect 1609 -94 1779 -34
rect 1925 -94 2095 -34
rect 2241 -94 2411 -34
rect 2557 -94 2727 -34
rect 2873 -94 3043 -34
rect 3189 -94 3249 -34
<< metal2 >>
rect 565 94 3503 114
rect 565 34 585 94
rect 3119 34 3503 94
rect 565 14 3503 34
rect 201 -16 3269 -14
rect 107 -34 3269 -16
rect 107 -36 455 -34
rect 107 -96 127 -36
rect 187 -94 455 -36
rect 515 -94 661 -34
rect 831 -94 977 -34
rect 1147 -94 1293 -34
rect 1463 -94 1609 -34
rect 1779 -94 1925 -34
rect 2095 -94 2241 -34
rect 2411 -94 2557 -34
rect 2727 -94 2873 -34
rect 3043 -94 3189 -34
rect 3249 -94 3269 -34
rect 187 -96 3269 -94
rect 107 -114 3269 -96
rect 107 -116 395 -114
rect -151 -812 -51 -792
rect -151 -872 -131 -812
rect -71 -872 -51 -812
rect -151 -892 -51 -872
rect 51 -812 151 -792
rect 51 -872 71 -812
rect 131 -872 151 -812
rect 51 -892 151 -872
<< labels >>
rlabel metal2 51 -892 151 -792 5 QN
rlabel metal2 -151 -892 -51 -792 5 Q
rlabel metal2 3403 14 3503 114 3 Vout
rlabel metal1 287 2336 387 2436 1 VDD
rlabel metal1 267 -1088 367 -988 5 VSS
<< end >>
