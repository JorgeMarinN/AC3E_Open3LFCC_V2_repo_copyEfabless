magic
tech sky130A
timestamp 1699136175
<< metal2 >>
rect 30400 100560 31270 100800
rect 31460 100560 32000 100800
rect 30400 98600 32000 100560
rect 32000 89060 33600 91800
rect 32240 88870 33600 89060
rect 32000 88000 33600 88870
rect 32000 34730 33600 35600
rect 32240 34540 33600 34730
rect 32000 31800 33600 34540
rect 31200 23438 32000 25400
rect 31451 23100 32000 23438
<< metal3 >>
rect 6000 128600 36000 131600
rect 0 99600 4000 126600
rect 33000 101600 36000 128600
rect 0 96800 30000 99600
rect 0 96600 31200 96800
rect 1000 95600 31200 96600
rect 1000 94800 31000 95600
rect 1000 93800 22000 94800
rect 0 90800 31200 93800
rect 0 63800 4200 90800
rect 33200 80000 36200 88800
rect 33200 61800 37200 80000
rect 6200 58800 37200 61800
rect 16000 58200 37200 58800
rect 16000 57600 37000 58200
rect 14800 57200 37000 57600
rect 16000 56600 37000 57200
rect 14800 53600 37200 56600
rect 8800 32800 12800 51600
rect 33600 34800 37200 53600
rect 8800 29800 31600 32800
rect 9000 28800 30000 29800
rect 9000 28400 31600 28800
rect 9000 27400 30000 28400
rect 8800 24400 30200 27400
rect 8800 5600 12400 24400
rect 33200 3600 36200 22400
rect 14400 600 36200 3600
<< metal4 >>
rect 6000 128600 36000 131600
rect 0 99600 4000 126600
rect 33000 101600 36000 128600
rect 0 96800 30000 99600
rect 0 96600 31200 96800
rect 1000 95600 31200 96600
rect 1000 94800 31000 95600
rect 1000 93800 22000 94800
rect 0 90800 31200 93800
rect 0 63800 4200 90800
rect 33200 80000 36200 88800
rect 33200 61800 37200 80000
rect 6200 58800 37200 61800
rect 16000 58200 37200 58800
rect 16000 57600 37000 58200
rect 14800 57200 37000 57600
rect 16000 56600 37000 57200
rect 14800 53600 37200 56600
rect 8800 32800 12800 51600
rect 33600 34800 37200 53600
rect 8800 29800 31600 32800
rect 9000 28800 30000 29800
rect 9000 28400 31600 28800
rect 9000 27400 30000 28400
rect 8800 24400 30200 27400
rect 8800 5600 12400 24400
rect 33200 3600 36200 22400
rect 14400 600 36200 3600
<< metal5 >>
rect 6000 128600 36000 131600
rect 0 99600 4000 126600
rect 33000 101600 36000 128600
rect 0 96800 30000 99600
rect 0 96600 31200 96800
rect 1000 95600 31200 96600
rect 1000 94800 31000 95600
rect 1000 93800 22000 94800
rect 0 90800 31200 93800
rect 0 63800 4200 90800
rect 33200 80000 36200 88800
rect 33200 61800 37200 80000
rect 6200 58800 37200 61800
rect 14000 58200 37200 58800
rect 14000 56600 37000 58200
rect 14000 56000 37200 56600
rect 14800 53600 37200 56000
rect 8800 32800 12800 51600
rect 33600 34800 37200 53600
rect 8800 29800 31600 32800
rect 9000 28800 30000 29800
rect 9000 28400 31600 28800
rect 9000 27400 30000 28400
rect 8800 24400 30200 27400
rect 8800 5600 12400 24400
rect 33200 3600 36200 22400
rect 14400 600 36200 3600
use nmos_waffle_32x32  nmos_waffle_32x32_0
timestamp 1698344533
transform 0 -1 31225 -1 0 22475
box -5925 -5975 22475 22425
use nmos_waffle_32x32  nmos_waffle_32x32_1
timestamp 1698344533
transform -1 0 31275 0 1 34775
box -5925 -5975 22475 22425
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1684343764
transform -1 0 31275 0 -1 88825
box -5925 -5975 31275 31225
use pmos_waffle_48x48  pmos_waffle_48x48_1
timestamp 1684343764
transform 0 -1 31225 1 0 101525
box -5925 -5975 31275 31225
<< labels >>
rlabel metal5 1000 94600 2000 95600 7 fc1
rlabel metal5 14800 56600 31200 57600 7 out
rlabel metal5 9800 28300 10800 29300 7 fc2
rlabel metal2 31200 24400 31700 25400 1 s4
rlabel metal5 34200 21400 35200 22400 1 VN
rlabel metal2 32600 31800 33600 32800 5 s3
rlabel metal2 32200 90800 33200 91800 1 s2
rlabel metal5 34000 101600 35000 102600 5 VP
rlabel metal2 31000 98600 32000 99600 5 s1
<< end >>
