magic
tech sky130A
magscale 1 2
timestamp 1699897858
<< checkpaint >>
rect -3932 125824 78332 269532
rect 0 97265 78332 125824
rect -22865 -5265 288465 97265
rect 92335 -22865 288465 -5265
<< obsactive >>
rect -18933 80852 284533 93333
rect -18933 74802 42950 80852
rect 51886 74802 62250 80852
rect 71186 74802 176150 80852
rect 185086 74802 196650 80852
rect 205586 74802 284533 80852
rect -18933 74400 284533 74802
rect -18933 17600 0 74400
rect 56800 17600 57600 74400
rect 114400 17600 115200 74400
rect -18933 0 115200 17600
rect 189600 0 191200 74400
rect 265600 0 284533 74400
rect -18933 -1333 284533 0
rect 96267 -18933 284533 -1333
<< metal1 >>
rect 2000 83200 212650 83800
rect 46450 83090 212650 83100
rect 46450 82910 46460 83090
rect 46640 82910 212650 83090
rect 46450 82900 212650 82910
rect 65750 82790 212650 82800
rect 65750 82610 65760 82790
rect 65940 82610 212650 82790
rect 65750 82600 212650 82610
rect 179650 82490 212650 82500
rect 179650 82310 179660 82490
rect 179840 82310 212650 82490
rect 179650 82300 212650 82310
rect 200150 82190 212650 82200
rect 200150 82010 200160 82190
rect 200340 82010 212650 82190
rect 200150 82000 212650 82010
rect 2000 81890 266550 81900
rect 2000 81410 46144 81890
rect 46210 81410 65444 81890
rect 65510 81410 179344 81890
rect 179410 81410 199844 81890
rect 199910 81410 266550 81890
rect 2000 81400 266550 81410
rect 2000 80700 212650 81300
<< via1 >>
rect 46460 82910 46640 83090
rect 65760 82610 65940 82790
rect 179660 82310 179840 82490
rect 200160 82010 200340 82190
rect 46144 81410 46210 81890
rect 65444 81410 65510 81890
rect 179344 81410 179410 81890
rect 199844 81410 199910 81890
rect 46144 79812 46210 80272
rect 47020 79612 47200 80192
rect 65444 79812 65510 80272
rect 66320 79612 66500 80192
rect 179344 79812 179410 80272
rect 180220 79612 180400 80192
rect 199844 79812 199910 80272
rect 200720 79612 200900 80192
<< metal2 >>
rect 5000 75990 6000 83800
rect 46450 83090 46650 83100
rect 46450 82910 46460 83090
rect 46640 82910 46650 83090
rect 46134 81890 46220 81900
rect 46134 81410 46144 81890
rect 46210 81410 46220 81890
rect 46134 80272 46220 81410
rect 46450 80532 46650 82910
rect 46134 79812 46144 80272
rect 46210 79812 46220 80272
rect 46134 79802 46220 79812
rect 47010 80192 47210 83800
rect 65750 82790 65950 82800
rect 65750 82610 65760 82790
rect 65940 82610 65950 82790
rect 47010 79612 47020 80192
rect 47200 79612 47210 80192
rect 65434 81890 65520 81900
rect 65434 81410 65444 81890
rect 65510 81410 65520 81890
rect 65434 80272 65520 81410
rect 65750 80532 65950 82610
rect 65434 79812 65444 80272
rect 65510 79812 65520 80272
rect 65434 79802 65520 79812
rect 66310 80192 66510 83800
rect 179650 82490 179850 82500
rect 179650 82310 179660 82490
rect 179840 82310 179850 82490
rect 47010 79602 47210 79612
rect 66310 79612 66320 80192
rect 66500 79612 66510 80192
rect 179334 81890 179420 81900
rect 179334 81410 179344 81890
rect 179410 81410 179420 81890
rect 179334 80272 179420 81410
rect 179650 80532 179850 82310
rect 179334 79812 179344 80272
rect 179410 79812 179420 80272
rect 179334 79802 179420 79812
rect 180210 80192 180410 83800
rect 200150 82190 200350 82200
rect 200150 82010 200160 82190
rect 200340 82010 200350 82190
rect 66310 79602 66510 79612
rect 180210 79612 180220 80192
rect 180400 79612 180410 80192
rect 199834 81890 199920 81900
rect 199834 81410 199844 81890
rect 199910 81410 199920 81890
rect 199834 80272 199920 81410
rect 200150 80532 200350 82010
rect 199834 79812 199844 80272
rect 199910 79812 199920 80272
rect 199834 79802 199920 79812
rect 200710 80192 200910 83800
rect 180210 79602 180410 79612
rect 200710 79612 200720 80192
rect 200900 79612 200910 80192
rect 200710 79602 200910 79612
rect 5000 75010 5010 75990
rect 5990 75010 6000 75990
rect 5000 75000 6000 75010
rect 260550 75990 261550 81900
rect 260550 75010 260560 75990
rect 261540 75010 261550 75990
rect 260550 75000 261550 75010
rect 47044 68772 47644 74902
rect 47044 68032 47074 68772
rect 47614 68032 47644 68772
rect 47044 63802 47644 68032
rect 66344 68772 66944 74902
rect 66344 68032 66374 68772
rect 66914 68032 66944 68772
rect 66344 66802 66944 68032
rect 180244 68772 180844 74902
rect 180244 68032 180274 68772
rect 180814 68032 180844 68772
rect 180244 66802 180844 68032
rect 200744 68772 201344 74902
rect 200744 68032 200774 68772
rect 201314 68032 201344 68772
rect 200744 63802 201344 68032
<< via2 >>
rect 5010 75010 5990 75990
rect 260560 75010 261540 75990
rect 47074 68032 47614 68772
rect 66374 68032 66914 68772
rect 180274 68032 180814 68772
rect 200774 68032 201314 68772
<< metal3 >>
rect 5000 75990 6000 76000
rect 5000 75010 5010 75990
rect 5990 75010 6000 75990
rect 5000 62000 6000 75010
rect 260550 75990 261550 76000
rect 260550 75010 260560 75990
rect 261540 75010 261550 75990
rect 47044 68772 47644 74902
rect 47044 68032 47074 68772
rect 47614 68032 47644 68772
rect 47044 63802 47644 68032
rect 66344 68772 66944 74902
rect 66344 68032 66374 68772
rect 66914 68032 66944 68772
rect 66344 66802 66944 68032
rect 180244 68772 180844 74902
rect 180244 68032 180274 68772
rect 180814 68032 180844 68772
rect 180244 66802 180844 68032
rect 200744 68772 201344 74902
rect 200744 68032 200774 68772
rect 201314 68032 201344 68772
rect 200744 63802 201344 68032
rect 260550 62000 261550 75010
<< via3 >>
rect 47074 68032 47614 68772
rect 66374 68032 66914 68772
rect 180274 68032 180814 68772
rect 200774 68032 201314 68772
<< metal4 >>
rect 47044 68772 47644 74902
rect 47044 68032 47074 68772
rect 47614 68032 47644 68772
rect 47044 63802 47644 68032
rect 66344 68772 66944 74902
rect 66344 68032 66374 68772
rect 66914 68032 66944 68772
rect 66344 66802 66944 68032
rect 180244 68772 180844 74902
rect 180244 68032 180274 68772
rect 180814 68032 180844 68772
rect 180244 66802 180844 68032
rect 200744 68772 201344 74902
rect 200744 68032 200774 68772
rect 201314 68032 201344 68772
rect 200744 63802 201344 68032
<< via4 >>
rect 47074 68032 47614 68772
rect 66374 68032 66914 68772
rect 180274 68032 180814 68772
rect 200774 68032 201314 68772
<< metal5 >>
rect 47044 68772 47644 74902
rect 47044 68032 47074 68772
rect 47614 68032 47644 68772
rect 47044 63802 47644 68032
rect 66344 68772 66944 74902
rect 66344 68032 66374 68772
rect 66914 68032 66944 68772
rect 66344 66802 66944 68032
rect 180244 68772 180844 74902
rect 180244 68032 180274 68772
rect 180814 68032 180844 68772
rect 180244 66802 180844 68032
rect 200744 68772 201344 74902
rect 200744 68032 200774 68772
rect 201314 68032 201344 68772
rect 200744 63802 201344 68032
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 196650 -1 0 80852
box 0 0 6050 8936
use level_shifter  level_shifter_1
timestamp 1666543010
transform 0 1 176150 -1 0 80852
box 0 0 6050 8936
use level_shifter  level_shifter_2
timestamp 1666543010
transform 0 1 62250 -1 0 80852
box 0 0 6050 8936
use level_shifter  level_shifter_3
timestamp 1666543010
transform 0 1 42950 -1 0 80852
box 0 0 6050 8936
use power_stage_1  power_stage_1_0
timestamp 1699136175
transform 0 1 0 1 0 0
box 0 0 74400 265600
<< labels >>
rlabel metal1 199450 80700 212650 81300 3 VLS
rlabel metal1 253350 81400 266550 81900 7 VDD
rlabel metal1 212450 82000 212650 82200 7 D1
rlabel metal1 212450 82300 212650 82500 7 D2
rlabel metal1 212450 82600 212650 82800 7 D3
rlabel metal1 212450 82900 212650 83100 7 D4
<< end >>
