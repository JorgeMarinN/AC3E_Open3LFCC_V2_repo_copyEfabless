
.subckt modulator CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT VGND
+ VPWR d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5]
.ends

