* NGSPICE file created from short_pulse_generator.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VPWR X VNB VPB
X0 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.33 as=0.213 ps=2.16 w=0.82 l=0.5
X1 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.217 pd=2.17 as=0.17 ps=1.36 w=0.82 l=0.5
X2 VPWR a_390_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.138 ps=1.27 w=1 l=0.15
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.36 as=0.27 ps=2.54 w=1 l=0.15
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.158 ps=1.33 w=1 l=0.15
X5 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=0.098 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.5
X6 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.01 as=0.113 ps=1.38 w=0.42 l=0.15
X7 VGND a_390_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.164 pd=1.62 as=0.0578 ps=0.695 w=0.42 l=0.15
X8 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=1.01 w=0.65 l=0.5
X9 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.098 ps=0.98 w=0.42 l=0.15
.ends

.subckt sp_delay sky130_fd_sc_hd__clkdlybuf4s50_2_0/A sky130_fd_sc_hd__clkdlybuf4s50_2_5/X
+ sky130_fd_sc_hd__tap_1_1/VPB VSUBS
Xsky130_fd_sc_hd__clkdlybuf4s50_2_0 sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_1/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_1 sky130_fd_sc_hd__clkdlybuf4s50_2_1/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_2/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_2 sky130_fd_sc_hd__clkdlybuf4s50_2_2/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_3/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_3 sky130_fd_sc_hd__clkdlybuf4s50_2_3/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_4/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_4 sky130_fd_sc_hd__clkdlybuf4s50_2_4/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_5/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_5 sky130_fd_sc_hd__clkdlybuf4s50_2_5/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_5/X VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
.ends

.subckt sp_delay2x VIN VOUT VSS VCC
Xsp_delay_0 VIN sp_delay_1/sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VCC VSS sp_delay
Xsp_delay_1 sp_delay_1/sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VOUT VCC VSS sp_delay
.ends

.subckt sp_delay_top VCC VIN VOUT VSS
Xsp_delay2x_0 VIN sp_delay2x_1/VIN VSS VCC sp_delay2x
Xsp_delay2x_1 sp_delay2x_1/VIN sp_delay2x_2/VIN VSS VCC sp_delay2x
Xsp_delay2x_2 sp_delay2x_2/VIN VOUT VSS VCC sp_delay2x
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VPWR X VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt short_pulse_generator VSS VCC Vin VFE VRE
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A VSS VCC sp_delay_top_0/VIN VSS
+ VCC sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_2_0 Vin VSS VCC sky130_fd_sc_hd__inv_2_0/Y VSS VCC sky130_fd_sc_hd__inv_2
Xsp_delay_top_0 VCC sp_delay_top_0/VIN sp_delay_top_0/VOUT VSS sp_delay_top
Xsky130_fd_sc_hd__and2_2_0 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_8_0/A VSS
+ VCC VRE VSS VCC sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__and2_2_1 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/A VSS
+ VCC VFE VSS VCC sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__inv_1_1 sp_delay_top_0/VOUT VSS VCC sky130_fd_sc_hd__inv_1_2/A VSS
+ VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_2_0/Y VSS VCC sky130_fd_sc_hd__inv_8_0/A
+ VSS VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VSS VCC sky130_fd_sc_hd__inv_1_2/Y
+ VSS VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_8_0/A VSS VCC sky130_fd_sc_hd__inv_1_3/Y
+ VSS VCC sky130_fd_sc_hd__inv_1
.ends

