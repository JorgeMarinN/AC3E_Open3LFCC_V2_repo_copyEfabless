magic
tech sky130A
timestamp 1698162338
<< obsactive >>
rect -9585 136794 46815 146794
rect -9585 100394 415 136794
rect 36815 100394 46815 136794
rect -9585 98794 46815 100394
rect -9585 62394 415 98794
rect 36815 62394 46815 98794
rect -9585 61194 46815 62394
rect -9585 31394 415 61194
rect 30215 52394 46815 61194
rect 30215 31394 40215 52394
rect -9585 30194 40215 31394
rect -9585 394 415 30194
rect 30215 394 40215 30194
rect -9585 -1000 40215 394
<< end >>
