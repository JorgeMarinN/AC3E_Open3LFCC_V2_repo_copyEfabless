* NGSPICE file created from power_stage_1.ext - technology: sky130A

.subckt pmos_source_in m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# m5_788_894# m4_0_0#
+ a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.86 ps=16.6 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=6.86 pd=16.6 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_drain_in m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.78 ps=18.8 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=2.78 pd=18.8 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_source_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.23 ps=16.3 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=6.23 pd=16.3 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_source_frame_lt m4_n1950_0# m4_648_1020# w_n1150_0# m5_n1950_0# m5_788_894#
+ m3_n1950_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_n1150_0# w_n1150_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=12.5 ps=32.6 w=4.38 l=0.5
.ends

.subckt pmos_drain_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# a_100_62#
+ m5_788_894# m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.03 ps=14.1 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.1 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_drain_frame_lt m4_648_1020# w_n1150_0# m3_n950_0# m4_n950_0# m5_n950_0#
+ m5_788_894# a_0_0# a_162_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_162_0# w_n1150_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=4.05 ps=28.2 w=4.38 l=0.5
.ends

.subckt pmos_waffle_48x48 a_n938_0# a_n1100_n1200# a_50762_0#
Xpmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_802 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_824 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_868 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_846 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_879 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_835 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_857 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_813 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_614 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_625 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_647 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_603 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_636 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_669 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_658 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_38 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1051 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1040 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_643 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_621 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_610 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_632 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_687 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_665 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_698 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_654 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_676 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_433 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_411 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_477 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_455 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_499 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_488 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_444 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_466 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_400 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_422 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_462 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_484 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_473 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_495 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_451 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_252 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_296 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_274 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_230 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_263 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_285 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_241 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_18 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_29 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_64 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_86 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_75 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_97 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_53 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1005 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1049 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1027 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1016 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1038 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_807 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_829 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_818 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_825 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_803 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_836 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_814 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_847 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_869 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_858 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_615 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_637 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_648 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_626 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_604 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_659 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1030 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1052 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_39 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1041 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_666 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_600 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_622 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_644 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_677 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_655 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_611 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_633 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_688 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_699 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_434 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_412 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_456 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_478 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_489 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_467 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_445 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_401 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_423 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_990 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_485 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_463 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_496 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_474 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_452 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_231 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_220 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_275 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_297 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_253 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_286 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_264 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_242 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_19 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_65 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_87 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_76 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_98 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_54 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1006 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1028 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1039 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1017 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_808 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_819 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_804 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_826 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_848 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_837 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_859 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_815 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_616 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_638 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_627 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_649 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_605 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1031 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1042 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1020 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1053 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_689 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_623 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_601 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_667 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_645 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_656 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_678 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_634 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_612 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_413 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_402 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_435 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_479 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_457 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_446 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_468 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_424 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_980 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_991 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_453 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_464 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_486 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_475 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_497 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_232 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_210 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_254 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_221 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_243 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_298 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_276 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_265 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_287 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_66 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_55 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_88 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_99 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_77 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1007 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1029 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1018 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_809 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_827 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_849 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_805 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_838 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_816 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_617 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_639 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_628 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_606 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1032 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1010 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1054 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1043 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1021 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_646 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_668 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_602 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_624 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_657 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_679 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_613 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_635 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_436 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_414 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_447 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_403 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_425 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_458 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_469 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_981 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_992 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_970 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_454 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_476 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_487 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_465 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_498 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_200 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_255 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_277 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_211 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_233 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_266 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_288 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_222 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_244 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_299 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_67 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_89 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_78 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_56 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1008 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1019 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_806 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_828 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_839 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_817 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_618 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_629 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_607 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1011 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1033 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1055 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1044 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1022 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1000 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_614 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_625 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_603 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_669 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_647 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_658 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_636 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_459 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_415 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_437 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_448 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_404 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_426 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_982 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_960 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_993 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_971 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_455 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_477 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_466 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_499 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_488 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_201 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_223 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_278 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_256 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_234 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_212 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_289 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_267 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_245 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_790 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_68 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_46 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_79 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_57 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1009 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_807 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_818 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_829 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_619 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_608 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1034 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1056 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1012 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1045 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1001 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1023 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_637 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_615 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_648 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_604 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_626 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_659 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_416 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_438 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_449 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_427 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_405 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_983 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_961 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_994 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_950 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_972 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_456 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_478 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_467 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_489 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_202 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_213 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_246 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_224 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_257 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_279 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_235 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_268 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_990 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_780 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_791 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_47 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_69 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_58 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_819 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_808 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_609 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1013 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1002 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1024 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1057 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1035 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1046 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_638 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_616 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_649 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_605 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_627 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_439 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_417 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_406 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_428 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_940 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_951 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_962 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_984 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_995 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_973 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_457 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_479 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_468 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_203 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_225 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_214 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_236 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_247 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_269 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_258 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_991 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_980 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_781 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_792 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_770 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_48 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_59 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_809 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1014 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1036 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1047 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1003 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1025 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_617 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_639 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_628 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_606 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_407 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_418 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_429 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_941 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_985 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_963 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_952 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_974 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_930 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_996 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_458 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_469 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_204 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_226 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_248 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_259 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_237 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_215 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_981 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_970 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_992 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_782 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_760 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_771 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_793 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_590 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_49 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1026 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1004 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1037 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1015 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1048 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_607 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_618 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_629 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_408 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_419 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_942 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_986 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_964 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_920 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_997 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_953 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_975 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_931 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_459 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_205 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_249 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_227 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_216 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_238 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_960 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_982 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_993 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_971 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_750 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_761 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_783 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_794 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_772 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_790 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_591 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_580 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1005 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1027 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1038 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1016 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1049 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_619 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_608 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_409 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_965 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_987 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_921 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_943 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_998 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_976 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_954 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_932 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_910 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_206 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_228 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_217 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_239 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_961 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_983 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_972 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_994 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_950 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_740 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_751 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_784 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_762 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_795 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_773 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_780 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_791 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_570 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_592 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_581 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1006 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1028 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1039 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1017 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_609 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_922 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_900 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_933 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_911 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_988 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_966 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_944 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_999 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_955 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_977 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_207 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_218 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_229 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_962 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_940 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_984 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_973 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_995 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_951 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_752 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_730 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_774 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_763 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_741 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_796 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_785 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_770 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_781 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_792 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_571 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_593 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_582 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_560 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_390 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1029 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1007 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1018 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_934 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_912 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_945 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_967 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_901 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_923 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_956 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_989 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_978 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_208 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_219 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_963 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_941 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_930 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_952 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_985 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_996 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_974 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_753 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_731 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_775 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_797 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_786 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_764 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_720 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_742 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_760 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_782 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_793 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_771 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_550 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_572 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_594 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_583 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_561 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_590 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_391 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_380 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1008 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1019 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_913 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_935 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_968 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_946 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_924 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_902 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_979 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_957 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_209 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_942 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_964 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_986 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_920 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_975 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_997 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_953 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_931 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_710 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_732 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_754 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_798 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_776 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_765 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_787 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_743 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_721 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_761 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_783 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_794 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_772 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_750 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_540 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_551 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_573 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_595 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_584 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_562 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_591 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_580 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_370 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_392 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_381 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1009 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_936 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_914 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_958 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_947 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_969 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_903 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_925 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_965 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_987 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_943 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_921 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_976 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_998 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_932 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_954 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_910 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_711 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_722 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_700 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_755 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_733 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_799 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_777 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_766 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_788 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_744 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_773 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_751 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_784 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_740 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_762 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_795 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_574 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_530 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_552 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_563 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_541 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_596 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_585 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_570 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_592 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_581 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_393 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_371 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_360 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_382 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_190 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_915 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_904 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_937 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_959 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_948 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_926 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_911 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_900 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_988 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_922 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_944 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_966 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_999 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_977 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_933 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_955 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_712 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_756 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_734 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_723 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_745 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_701 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_778 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_789 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_767 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_730 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_752 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_741 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_774 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_785 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_763 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_796 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_597 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_531 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_553 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_575 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_586 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_542 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_564 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_520 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_571 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_593 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_582 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_560 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_361 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_394 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_372 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_350 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_383 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_180 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_191 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_916 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_938 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_949 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_927 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_905 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_912 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_945 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_923 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_901 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_934 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_989 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_967 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_978 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_956 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_735 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_757 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_779 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_713 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_768 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_746 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_724 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_702 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_731 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_775 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_753 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_786 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_742 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_764 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_720 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_797 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_554 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_532 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_598 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_576 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_510 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_587 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_565 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_543 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_521 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_550 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_594 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_572 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_583 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_561 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_340 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_384 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_362 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_395 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_351 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_373 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_181 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_170 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_192 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_939 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_917 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_906 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_928 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_913 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_957 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_935 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_968 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_924 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_946 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_902 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_979 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_758 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_736 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_714 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_769 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_725 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_747 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_703 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_732 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_710 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_776 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_754 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_798 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_787 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_743 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_765 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_721 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_522 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_500 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_511 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_577 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_599 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_555 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_533 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_588 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_566 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_544 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_551 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_573 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_595 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_562 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_584 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_540 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_341 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_363 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_352 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_374 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_330 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_385 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_396 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_160 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_182 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_171 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_193 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_918 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_907 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_929 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_914 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_936 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_958 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_969 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_947 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_925 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_903 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_704 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_715 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_737 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_759 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_726 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_748 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_711 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_700 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_733 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_755 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_777 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_799 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_788 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_766 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_744 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_722 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_523 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_501 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_545 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_556 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_534 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_512 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_578 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_589 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_567 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_530 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_552 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_541 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_574 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_596 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_585 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_563 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_342 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_320 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_364 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_386 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_397 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_375 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_353 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_331 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_183 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_161 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_194 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_172 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_150 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_919 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_908 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_915 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_959 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_937 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_926 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_948 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_904 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_738 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_716 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_727 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_705 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_749 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_712 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_734 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_723 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_701 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_778 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_756 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_789 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_745 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_767 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_502 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_524 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_546 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_568 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_579 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_557 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_535 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_513 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_531 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_553 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_575 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_586 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_564 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_542 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_520 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_597 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_321 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_343 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_387 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_365 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_398 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_354 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_376 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_332 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_310 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_140 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_184 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_162 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_173 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_195 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_151 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_909 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_916 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_927 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_905 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_938 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_949 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_706 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_717 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_739 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_728 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_735 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_757 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_713 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_746 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_768 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_702 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_724 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_779 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_525 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_503 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_547 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_569 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_536 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_558 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_514 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_554 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_576 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_598 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_532 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_510 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_565 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_587 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_543 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_521 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_322 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_300 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_311 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_344 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_388 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_366 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_399 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_355 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_377 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_333 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_163 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_141 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_130 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_152 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_185 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_196 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_174 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_917 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_939 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_928 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_906 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_707 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_729 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_718 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_758 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_714 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_736 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_769 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_747 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_703 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_725 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_504 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_526 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_548 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_559 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_537 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_515 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_500 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_522 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_577 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_555 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_599 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_533 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_511 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_588 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_566 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_544 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_301 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_323 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_345 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_356 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_334 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_312 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_367 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_389 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_378 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_890 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_131 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_186 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_164 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_142 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_120 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_197 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_175 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_153 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_918 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_929 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_907 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_708 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_719 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_715 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_759 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_737 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_748 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_726 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_704 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_505 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_527 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_538 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_516 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_549 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_501 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_523 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_534 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_512 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_545 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_578 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_556 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_589 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_567 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_324 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_302 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_368 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_346 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_357 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_379 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_335 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_313 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_891 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_880 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_110 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_154 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_132 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_165 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_187 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_121 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_143 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_176 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_198 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_919 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_908 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_709 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_716 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_705 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_738 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_749 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_727 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_528 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_506 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_539 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_517 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_502 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_524 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_546 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_568 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_557 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_535 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_513 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_579 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_347 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_369 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_303 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_325 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_358 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_314 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_336 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_870 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_892 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_881 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_111 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_122 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_100 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_155 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_133 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_177 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_188 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_166 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_144 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_199 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_909 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_706 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_728 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_739 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_717 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_507 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_529 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_518 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_503 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_525 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_547 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_569 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_558 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_536 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_514 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_304 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_315 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_348 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_326 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_359 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_337 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_860 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_893 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_871 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_882 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_112 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_134 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_145 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_123 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_101 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_156 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_178 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_167 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_189 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_690 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_0 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_729 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_707 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_718 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_508 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_519 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_504 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_526 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_548 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_559 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_537 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_515 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_338 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_316 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_305 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_327 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_349 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_850 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_872 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_861 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_883 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_894 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_113 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_157 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_135 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_179 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_168 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_124 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_146 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_102 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_890 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_691 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_680 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_lt_1 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_40 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_708 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_719 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_509 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_505 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_516 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_527 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_549 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_538 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_339 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_317 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_306 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_328 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_873 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_895 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_851 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_884 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_862 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_840 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_114 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_158 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_136 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_169 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_125 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_147 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_103 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_891 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_880 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_692 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_670 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_681 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_2 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_30 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_41 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_709 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_528 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_506 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_539 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_517 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_318 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_329 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_307 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1050 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_896 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_830 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_874 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_852 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_863 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_885 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_841 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_104 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_137 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_159 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_115 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_148 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_126 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_870 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_892 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_881 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_660 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_671 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_693 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_682 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_40 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_3 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_490 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_42 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_20 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_31 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_507 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_529 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_518 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_319 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1051 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1040 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_308 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_842 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_820 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_831 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_853 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_875 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_897 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_864 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_886 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_116 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_127 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_105 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_138 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_149 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_871 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_893 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_882 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_860 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_661 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_683 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_672 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_650 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_694 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_41 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_4 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_690 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_480 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_491 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_32 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_10 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_43 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_21 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_508 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_519 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_309 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1052 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1030 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1041 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_821 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_843 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_854 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_832 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_810 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_865 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_876 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_898 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_887 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_117 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_139 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_128 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_106 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_850 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_872 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_861 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_894 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_883 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_640 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_662 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_684 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_673 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_695 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_651 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_42 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_5 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_691 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_680 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_481 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_492 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_470 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_22 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_33 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_11 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_44 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_90 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_509 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1031 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1053 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1042 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1020 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_800 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_844 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_822 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_888 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_866 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_899 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_855 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_877 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_811 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_833 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_118 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_129 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_107 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_873 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_895 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_851 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_884 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_840 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_862 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_663 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_641 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_685 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_674 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_696 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_630 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_652 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_43 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_6 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_692 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_670 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_681 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_482 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_460 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_493 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_471 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_290 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_34 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_12 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_45 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_23 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_91 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_80 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1010 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1054 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1032 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1021 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1043 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_801 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_845 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_823 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_867 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_889 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_878 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_856 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_812 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_834 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_108 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_119 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_896 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_830 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_852 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_874 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_885 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_863 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_841 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_620 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_631 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_664 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_642 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_686 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_697 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_675 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_653 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_44 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_7 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_660 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_693 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_671 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_682 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_461 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_483 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_472 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_450 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_494 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_490 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_280 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_291 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_24 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_35 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_13 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_92 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_70 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_81 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1011 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1033 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1022 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1000 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1055 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1044 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_802 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_824 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_813 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_846 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_868 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_857 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_879 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_835 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_109 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_820 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_853 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_831 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_897 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_875 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_886 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_864 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_842 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_643 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_665 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_621 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_654 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_632 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_610 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_687 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_676 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_698 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_34 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_45 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_8 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_661 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_650 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_683 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_694 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_672 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_462 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_440 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_484 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_495 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_473 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_451 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_480 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_491 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_292 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_270 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_281 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_36 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_14 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_25 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_71 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_93 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_82 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_60 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1034 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1056 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1012 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1045 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1023 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1001 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_803 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_847 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_825 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_814 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_836 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_869 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_858 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_821 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_843 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_832 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_854 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_810 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_865 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_876 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_898 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_887 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_666 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_688 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_600 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_644 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_622 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_677 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_699 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_633 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_655 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_611 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_35 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_9 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_640 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_684 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_662 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_695 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_651 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_673 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_430 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_485 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_441 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_463 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_496 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_452 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_474 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_481 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_470 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_492 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_293 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_271 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_15 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_260 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_282 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_26 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_37 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_50 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_94 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_72 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_83 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_61 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1057 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1035 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1013 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1024 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1046 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1002 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_804 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_848 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_826 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_859 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_815 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_837 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_822 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_800 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_844 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_866 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_877 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_855 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_833 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_811 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_899 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_888 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_689 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_623 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_645 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_667 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_601 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_678 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_634 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_656 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_612 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_36 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_641 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_663 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_685 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_696 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_674 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_652 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_630 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_431 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_420 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_453 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_486 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_464 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_442 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_497 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_475 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_482 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_460 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_493 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_471 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_250 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_272 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_283 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_261 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_38 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_16 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_294 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_27 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_62 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_73 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_51 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_84 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_95 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1003 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1014 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1036 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1047 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1025 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_827 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_849 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_805 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_838 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_816 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_801 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_823 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_867 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_845 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_889 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_878 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_834 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_856 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_812 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_602 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_613 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_646 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_624 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_668 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_679 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_657 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_635 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1050 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_37 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_620 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_642 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_686 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_664 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_697 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_653 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_675 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_631 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_410 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_432 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_454 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_443 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_465 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_421 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_476 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_487 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_498 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_461 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_450 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_483 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_472 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_494 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_251 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_295 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_273 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_262 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_284 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_240 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_28 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_39 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_17 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_63 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_85 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_96 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_74 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_52 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1004 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1015 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1037 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1048 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1026 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_806 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_828 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_817 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_839 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
X0 a_50762_0# a_n1100_n1200# a_n938_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X1 a_n938_0# a_n1100_n1200# a_50762_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_50762_0# a_n1100_n1200# a_n938_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_50762_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt nmos_source_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.86 ps=16.6 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=6.86 pd=16.6 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_drain_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# a_100_62#
+ m5_788_894# m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.78 ps=18.8 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.78 pd=18.8 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020# a_1550_0#
X0 a_162_1100# a_0_0# a_100_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.03 ps=14.1 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.1 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_lt m4_n1950_0# m4_648_1020# m5_n1950_0# a_n950_0# m5_788_894#
+ m3_n1950_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_n950_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=12.5 ps=32.6 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.23 ps=16.3 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=6.23 pd=16.3 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_lt m4_648_1020# m3_n950_0# a_n950_0# m4_n950_0# m5_n950_0#
+ m5_788_894# a_0_0# a_162_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_162_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=4.05 ps=28.2 w=4.38 l=0.5
.ends

.subckt nmos_waffle_32x32 a_33162_0# a_n938_0# a_n1100_n1200#
Xnmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_371 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_382 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_360 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_393 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_190 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_372 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_383 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_350 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_361 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_394 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_191 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_180 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_373 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_340 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_384 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_395 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_351 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_362 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_192 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_170 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_181 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_374 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_341 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_385 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_396 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_352 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_330 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_363 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_193 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_160 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_171 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_182 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_342 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_386 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_353 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_397 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_320 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_375 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_331 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_364 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_161 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_172 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_150 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_183 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_194 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_0 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_343 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_387 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_310 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_398 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_354 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_365 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_321 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_376 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_332 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_20 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_162 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_173 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_195 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_151 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_184 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_140 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_344 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_388 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_311 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_399 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_355 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_366 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_322 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_300 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_1 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_377 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_333 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_10 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_163 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_130 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_21 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_174 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_185 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_196 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_152 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_141 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_389 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_312 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_356 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_323 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_367 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_345 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_2 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_301 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_378 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_334 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_22 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_164 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_131 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_175 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_186 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_142 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_120 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_197 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_153 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_11 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_313 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_3 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_302 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_357 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_368 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_324 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_335 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_346 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_379 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_12 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_132 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_176 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_23 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_143 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_187 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_121 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_165 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_198 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_154 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_110 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_4 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_314 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_358 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_369 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_325 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_336 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_347 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_303 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_24 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_133 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_177 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_100 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_188 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_144 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_13 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_166 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_122 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_111 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_155 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_199 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_5 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_359 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_326 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_337 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_315 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_348 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_304 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_14 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_134 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_178 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_25 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_101 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_189 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_145 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_156 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_112 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_167 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_123 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_327 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_338 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_305 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_6 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_0 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_316 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_349 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_26 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_179 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_102 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_146 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_113 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_157 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_15 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_135 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_168 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_124 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_1 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_328 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_339 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_306 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_317 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_7 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_frame_lt_16 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_103 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_27 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_147 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_158 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_114 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_136 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_169 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_125 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_90 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_329 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_307 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_2 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_8 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_318 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_28 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_104 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_148 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_159 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_115 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_17 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_126 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_137 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_0 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_91 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_80 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_9 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_3 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_308 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_319 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_18 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_29 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_149 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_116 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_127 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_105 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_138 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_1 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_70 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_92 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_81 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_309 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_4 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_117 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_19 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_128 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_106 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_139 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_2 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_71 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_82 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_60 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_93 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_5 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_118 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_129 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_107 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_3 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_290 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_72 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_83 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_61 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_94 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_50 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_6 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_119 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_108 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_4 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_280 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_291 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_73 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_40 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_84 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_62 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_51 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_95 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_7 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_109 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_440 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_5 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_281 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_292 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_270 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_74 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_41 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_85 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_96 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_52 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_30 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_63 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_8 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_430 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_441 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_6 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_282 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_293 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_260 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_271 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_42 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_86 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_53 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_97 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_31 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_75 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_64 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_20 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_9 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_431 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_442 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_420 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_7 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_283 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_250 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_294 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_261 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_272 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_43 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_87 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_10 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_98 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_54 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_76 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_32 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_21 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_65 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_432 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_443 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_410 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_421 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_8 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_284 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_251 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_295 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_262 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_240 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_273 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_44 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_11 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_55 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_22 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_33 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_88 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_99 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_66 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_77 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_20 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_400 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_411 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_422 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_433 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_444 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_9 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_252 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_296 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_263 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_230 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_285 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_241 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_274 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_89 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_12 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_56 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_23 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_67 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_45 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_78 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_34 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_21 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_10 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_434 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_401 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_445 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_412 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_423 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_253 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_297 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_220 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_264 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_275 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_231 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_286 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_242 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_20 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_13 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_57 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_68 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_24 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_46 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_79 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_35 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_11 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_22 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_0 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_402 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_446 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_413 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_435 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_424 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_254 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_298 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_221 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_21 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_265 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_276 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_232 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_10 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_210 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_287 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_243 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_14 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_58 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_69 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_25 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_36 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_47 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_23 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_1 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_12 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_403 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_447 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_414 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_425 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_436 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_299 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_222 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_266 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_233 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_277 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_200 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_255 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_211 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_288 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_244 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_59 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_26 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_37 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_11 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_22 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_15 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_48 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_13 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_2 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_lt_24 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_404 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_448 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_415 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_426 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_437 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_223 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_267 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_278 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_234 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_245 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_201 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_256 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_212 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_289 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_23 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_27 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_38 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_16 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_12 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_49 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_25 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_14 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_3 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_416 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_427 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_405 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_438 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_449 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_224 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_268 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_279 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_235 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_246 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_202 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_257 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_213 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_13 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_24 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_28 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_39 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_17 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_15 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_26 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_4 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_417 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_428 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_406 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_439 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_269 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_236 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_203 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_247 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_225 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_258 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_214 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_25 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_14 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_29 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_18 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_27 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_16 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_5 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_418 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_429 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_407 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_204 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_237 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_248 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_15 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_215 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_26 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_226 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_259 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_19 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_17 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_6 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_lt_28 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_419 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_408 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_238 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_249 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_205 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_216 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_227 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_27 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_16 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_29 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_18 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_7 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_409 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_239 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_206 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_217 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_228 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_17 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_28 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_19 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_8 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_207 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_218 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_229 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_29 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_18 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_390 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_9 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_208 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_219 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_19 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_380 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_391 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_209 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_370 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_381 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_392 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
X0 a_n938_0# a_n1100_n1200# a_33162_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X1 a_33162_0# a_n1100_n1200# a_n938_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_33162_0# a_n1100_n1200# a_n938_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_33162_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt power_stage_1
Xpmos_waffle_48x48_0 out s2 fc1 pmos_waffle_48x48
Xpmos_waffle_48x48_1 fc1 s1 VP pmos_waffle_48x48
Xnmos_waffle_32x32_0 VN fc2 s4 nmos_waffle_32x32
Xnmos_waffle_32x32_1 fc2 out s3 nmos_waffle_32x32
.ends

