* NGSPICE file created from Modulator.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_2 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.223 pd=2.21 as=0.121 ps=1.16 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.121 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VPB VNB VGND VPWR
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 VNB VPB VGND VPWR A1 A0 S0 A3 A2 S1 X
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0852 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.269 pd=2.12 as=0.0921 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0921 pd=0.99 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0852 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0901 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0901 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.151 ps=1.28 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151 pd=1.28 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.5 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.169 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.168 ps=1.5 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.5 as=0.109 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_2 VPB VNB VGND VPWR Y A B_N
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR VNB VPB A X B_N
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.266 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 VPB VNB A1 A2 A3 Y B1 VPWR VGND
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VPB VNB VGND VPWR A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.263 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.213 ps=1.42 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 VPB VNB VGND VPWR C_N B Y A
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_2 VPB VNB VGND VPWR A1 A2 Y B2 B1
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VNB VPB VGND VPWR A2 A1 B1 B2 Y C1
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_4 VNB VPB VGND VPWR B1_N A2 X A1
X0 a_1021_47# A1 a_205_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND A2 a_1021_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND a_42_47# a_205_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_861_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.101 ps=0.96 w=0.65 l=0.15
X7 a_205_21# A1 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0747 ps=0.88 w=0.65 l=0.15
X8 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_603_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND B1_N a_42_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.25 ps=2.07 w=0.65 l=0.15
X11 VPWR A2 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_603_297# a_42_47# a_205_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X14 a_205_21# a_42_47# a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.263 pd=1.46 as=0.091 ps=0.93 w=0.65 l=0.15
X16 VPWR B1_N a_42_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X17 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR A1 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_603_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_205_21# a_42_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.263 ps=1.46 w=0.65 l=0.15
X21 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_2 VNB VPB VGND VPWR B1 B2 A3 A2 A1 X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.14 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.123 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 VNB VPB VGND VPWR X B1 A2 A1 A3
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.1 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0536 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VPB VNB VGND VPWR Y B C A_N
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125 ps=1.03 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 VPB VNB VGND VPWR X B1 A4 A3 A2 A1
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.123 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.127 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VPB VNB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VNB VPB VPWR VGND X S A1 A0
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.109 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.275 ps=1.5 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_1 VNB VPB VGND VPWR A1 A2 A3 A4 Y B1
X0 a_348_297# A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.312 ps=1.62 w=1 l=0.15
X1 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.114 ps=1 w=0.65 l=0.15
X2 a_193_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A1 a_432_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.175 ps=1.35 w=1 l=0.15
X4 VGND A4 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.203 ps=1.27 w=0.65 l=0.15
X5 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_432_297# A2 a_348_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 VPWR VGND VPB VNB X A
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt Modulator CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT VGND
+ VPWR d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5]
XFILLER_0_27_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1270_ VGND VPWR _0180_ _0629_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0985_ VPWR VGND VPWR VGND _0058_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ VGND VPWR _0285_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ _0284_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1322_ VPWR VGND VPWR VGND Signal_Generator_1_270phase_inst.count\[5\] _0105_ _0019_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1253_ VPWR VGND VPWR VGND _0455_ _0454_ Dead_Time_Generator_inst_4.count_dt\[0\]
+ _0617_ sky130_fd_sc_hd__a21oi_1
X_1184_ VPWR VGND VGND VPWR _0563_ _0565_ _0564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0968_ VPWR VGND VGND VPWR Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\]
+ _0430_ sky130_fd_sc_hd__nor2_1
X_0899_ VPWR VGND VPWR VGND _0381_ _0367_ _0378_ _0038_ Signal_Generator_2_180phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0822_ VPWR VGND VPWR VGND Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[2\]
+ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[0\]
+ _0323_ sky130_fd_sc_hd__or4_2
XFILLER_0_28_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ VPWR VGND VPWR VGND _0271_ _0262_ _0269_ _0023_ Signal_Generator_1_90phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0684_ VGND VPWR _0143_ _0221_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1305_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0088_ net49
+ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
XFILLER_0_36_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1236_ VPWR VGND _0606_ _0604_ _0603_ VPWR VGND sky130_fd_sc_hd__and2_1
X_1098_ VPWR VGND VPWR VGND _0114_ _0499_ sky130_fd_sc_hd__inv_2
X_1167_ VPWR VGND _0549_ _0548_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ _0460_ Shift_Register_Inst.data_out\[8\] Shift_Register_Inst.data_out\[7\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0805_ VPWR VGND VPWR VGND _0310_ _0304_ _0309_ _0015_ Signal_Generator_1_270phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0736_ _0259_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0239_ Signal_Generator_1_0phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_0667_ VGND VPWR VPWR VGND _0190_ _0196_ Shift_Register_Inst.shift_state\[1\] _0209_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1219_ VPWR VGND VPWR VGND _0585_ Dead_Time_Generator_inst_2.count_dt\[3\] Dead_Time_Generator_inst_2.count_dt\[4\]
+ _0591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold41 net66 Signal_Generator_2_180phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net77 Signal_Generator_2_90phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 net55 Dead_Time_Generator_inst_1.count_dt\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1004_ VPWR VGND _0445_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_44_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0719_ VPWR VGND VGND VPWR _0246_ _0245_ _0242_ sky130_fd_sc_hd__or2_1
Xoutput20 VGND VPWR net20 PMOS1_PS1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0984_ VPWR VGND VPWR VGND _0057_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_142 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1321_ VGND VPWR VPWR VGND clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0018_
+ _0104_ Signal_Generator_1_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1252_ VGND VPWR _0616_ _0454_ Dead_Time_Generator_inst_4.count_dt\[0\] _0455_ VPWR
+ VGND sky130_fd_sc_hd__and3_1
X_1183_ VPWR VGND VGND VPWR _0564_ Dead_Time_Generator_inst_1.count_dt\[1\] net32
+ sky130_fd_sc_hd__or2_1
XFILLER_0_24_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0967_ VGND VPWR VGND VPWR net20 net22 _0428_ net17 net15 Shift_Register_Inst.data_out\[9\]
+ _0429_ sky130_fd_sc_hd__mux4_1
X_0898_ VPWR VGND VPWR VGND _0380_ _0379_ _0370_ _0381_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0752_ VPWR VGND VGND VPWR _0271_ net35 _0270_ sky130_fd_sc_hd__or2_1
X_0821_ VPWR VGND _0019_ _0306_ Signal_Generator_1_270phase_inst.direction Signal_Generator_1_270phase_inst.count\[4\]
+ _0322_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ VGND VPWR VPWR VGND _0221_ Shift_Register_Inst.data_out\[9\] _0220_ _0182_
+ sky130_fd_sc_hd__mux2_1
X_1304_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[1\] _0087_ _0022_
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1166_ VPWR VGND VPWR VGND _0542_ _0547_ _0548_ _0514_ net45 sky130_fd_sc_hd__or4b_2
X_1235_ VGND VPWR _0605_ _0603_ Dead_Time_Generator_inst_3.count_dt\[0\] _0604_ VPWR
+ VGND sky130_fd_sc_hd__and3_1
X_1097_ VPWR VGND VPWR VGND _0113_ _0499_ sky130_fd_sc_hd__inv_2
X_1020_ VPWR VGND VGND VPWR _0459_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\]
+ sky130_fd_sc_hd__nor2b_2
XPHY_EDGE_ROW_28_Left_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0735_ VGND VPWR VPWR VGND _0004_ _0257_ _0256_ Signal_Generator_1_0phase_inst.direction
+ _0241_ _0258_ sky130_fd_sc_hd__a32o_1
X_0804_ VGND VPWR VGND VPWR _0307_ _0310_ _0309_ sky130_fd_sc_hd__or2b_1
X_0666_ VGND VPWR Shift_Register_Inst.data_out\[5\] _0208_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_1218_ VGND VPWR _0167_ _0590_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1149_ VPWR VGND VGND VPWR _0530_ _0512_ _0511_ _0514_ _0531_ sky130_fd_sc_hd__o22a_1
Xhold31 net56 Signal_Generator_2_270phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 net78 Signal_Generator_1_0phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net45 _0546_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 net67 Dead_Time_Generator_inst_1.dt\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ VPWR VGND VPWR VGND _0075_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0718_ VPWR VGND VGND VPWR Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ _0245_ sky130_fd_sc_hd__nor2_1
X_0649_ VPWR VGND _0197_ _0196_ Shift_Register_Inst.shift_state\[0\] VPWR VGND sky130_fd_sc_hd__and2_1
Xoutput21 VGND VPWR net21 PMOS1_PS2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0983_ VPWR VGND VPWR VGND _0056_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1320_ VGND VPWR VPWR VGND clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0017_
+ _0103_ Signal_Generator_1_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1182_ VPWR VGND VGND VPWR Dead_Time_Generator_inst_1.count_dt\[1\] _0563_ net32
+ sky130_fd_sc_hd__nand2_1
X_1251_ VGND VPWR _0175_ _0615_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0897_ VPWR VGND _0380_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[1\]
+ net65 Signal_Generator_2_180phase_inst.count\[3\] VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_40_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0966_ VPWR VGND VPWR VGND _0428_ Shift_Register_Inst.data_out\[10\] sky130_fd_sc_hd__inv_2
XFILLER_0_10_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0751_ VGND VPWR VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0270_ _0263_
+ sky130_fd_sc_hd__xor2_1
X_0820_ _0322_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0302_ Signal_Generator_1_270phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_1303_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[0\] _0086_ _0021_
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_0682_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[2\] _0209_ _0188_ _0220_
+ sky130_fd_sc_hd__or3_1
X_1096_ VPWR VGND VPWR VGND _0112_ _0499_ sky130_fd_sc_hd__inv_2
X_1165_ VGND VPWR _0547_ _0521_ _0529_ _0528_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1234_ VGND VPWR VGND VPWR net30 _0604_ Dead_Time_Generator_inst_3.count_dt\[4\]
+ sky130_fd_sc_hd__or2b_1
X_0949_ VPWR VGND _0417_ _0416_ _0410_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_33_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0734_ VGND VPWR _0239_ _0258_ Signal_Generator_1_0phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_0803_ VPWR VGND VGND VPWR _0309_ _0308_ _0305_ sky130_fd_sc_hd__or2_1
X_0665_ VGND VPWR _0148_ _0207_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_74 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1079_ VPWR VGND VPWR VGND _0096_ _0498_ sky130_fd_sc_hd__inv_2
X_1217_ VGND VPWR _0590_ _0549_ _0545_ _0589_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1148_ VPWR VGND VPWR VGND _0529_ _0530_ _0521_ _0528_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_45_Left_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold43 net68 Dead_Time_Generator_inst_3.count_dt\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net35 _0265_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net57 Signal_Generator_1_180phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net46 _0548_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net79 Shift_Register_Inst.shift_state\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1002_ VPWR VGND VPWR VGND _0074_ _0444_ sky130_fd_sc_hd__inv_2
X_0717_ VPWR VGND VPWR VGND _0000_ net60 sky130_fd_sc_hd__inv_2
X_0648_ VGND VPWR _0185_ net72 _0196_ Shift_Register_Inst.shift_state\[1\] VPWR VGND
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 VGND VPWR net22 PMOS2_PS1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0982_ VPWR VGND _0443_ _0442_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_22_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1250_ VGND VPWR _0615_ _0548_ _0544_ _0614_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1181_ VPWR VGND VPWR VGND _0158_ _0562_ net32 _0545_ _0549_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_24_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0896_ VPWR VGND VPWR VGND _0379_ _0369_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ VPWR VGND VPWR VGND _0427_ Shift_Register_Inst.data_out\[12\] sky130_fd_sc_hd__inv_2
XFILLER_0_10_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0750_ VGND VPWR VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] _0269_ net48
+ sky130_fd_sc_hd__xor2_1
X_0681_ VGND VPWR _0144_ _0219_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1302_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.direction _0085_ net36
+ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
X_1233_ VPWR VGND VPWR VGND _0595_ net38 _0603_ _0600_ _0601_ _0602_ sky130_fd_sc_hd__a221o_1
X_1164_ VGND VPWR _0546_ _0526_ _0522_ _0527_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1095_ VPWR VGND VPWR VGND _0111_ _0499_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0948_ VGND VPWR VPWR VGND _0416_ net3 Shift_Register_Inst.data_out\[13\] Dead_Time_Generator_inst_2.go
+ sky130_fd_sc_hd__mux2_1
X_0879_ VPWR VGND VPWR VGND _0366_ Signal_Generator_2_180phase_inst.direction sky130_fd_sc_hd__inv_2
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0802_ VPWR VGND VGND VPWR Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ _0308_ sky130_fd_sc_hd__nor2_1
X_0733_ VPWR VGND VGND VPWR _0257_ Signal_Generator_1_0phase_inst.count\[4\] _0243_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0664_ VGND VPWR VPWR VGND _0207_ Dead_Time_Generator_inst_1.dt\[4\] _0206_ _0182_
+ sky130_fd_sc_hd__mux2_1
X_1216_ VGND VPWR _0585_ _0589_ _0569_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_1078_ VPWR VGND _0498_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
X_1147_ VPWR VGND VGND VPWR _0519_ _0529_ _0520_ sky130_fd_sc_hd__nand2_1
Xhold22 net47 Signal_Generator_1_90phase_inst.count\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net36 _0027_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold44 net69 _0173_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 net80 Signal_Generator_1_270phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 net58 Signal_Generator_1_270phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1001_ VPWR VGND VPWR VGND _0073_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0716_ VPWR VGND VGND VPWR _0241_ _0244_ _0006_ sky130_fd_sc_hd__nor2_1
X_0647_ VPWR VGND VGND VPWR _0192_ _0195_ _0154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput23 VGND VPWR net23 PMOS2_PS2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0981_ VPWR VGND _0442_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1180_ VPWR VGND VGND VPWR Dead_Time_Generator_inst_1.count_dt\[0\] _0561_ _0562_
+ sky130_fd_sc_hd__nor2_1
X_0964_ VGND VPWR net20 _0426_ VPWR VGND sky130_fd_sc_hd__buf_1
X_0895_ VPWR VGND VGND VPWR _0365_ _0378_ _0377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0680_ VGND VPWR VPWR VGND _0219_ _0217_ _0218_ _0182_ sky130_fd_sc_hd__mux2_1
X_1301_ VGND VPWR VPWR VGND clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0005_
+ _0084_ Signal_Generator_1_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_2
X_1232_ _0602_ Dead_Time_Generator_inst_3.count_dt\[4\] net64 VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and2b_1
X_1094_ VPWR VGND VPWR VGND _0110_ _0499_ sky130_fd_sc_hd__inv_2
X_1163_ VPWR VGND _0545_ _0544_ VPWR VGND sky130_fd_sc_hd__buf_2
X_0947_ VGND VPWR net23 _0415_ VPWR VGND sky130_fd_sc_hd__buf_1
X_0878_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[2\]
+ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[0\]
+ _0365_ sky130_fd_sc_hd__or4_2
X_0801_ VPWR VGND VPWR VGND _0014_ net58 sky130_fd_sc_hd__inv_2
XFILLER_0_21_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0732_ VGND VPWR VPWR VGND Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0253_ _0256_ sky130_fd_sc_hd__or3b_1
X_0663_ VPWR VGND VPWR VGND _0184_ _0193_ _0183_ _0206_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ VGND VPWR _0166_ _0588_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1146_ VPWR VGND VPWR VGND _0526_ _0522_ _0527_ _0528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1077_ VPWR VGND VPWR VGND _0095_ _0497_ sky130_fd_sc_hd__inv_2
Xhold12 net37 RST VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net48 _0266_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 net70 Signal_Generator_1_180phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 net59 Dead_Time_Generator_inst_3.count_dt\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ VPWR VGND VPWR VGND _0072_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0715_ VGND VPWR _0244_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.count\[5\]
+ _0243_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0646_ VPWR VGND _0195_ _0191_ _0189_ VPWR VGND sky130_fd_sc_hd__and2_1
X_1129_ VPWR VGND VPWR VGND _0511_ _0510_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 VGND VPWR net24 PMOS_PS3 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0980_ VGND VPWR net2 _0441_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_274 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR net26 clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_19_Left_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0894_ VPWR VGND net65 Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[2\]
+ _0377_ Signal_Generator_2_180phase_inst.count\[3\] VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0963_ VPWR VGND VGND VPWR _0426_ _0419_ _0423_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1300_ VGND VPWR VPWR VGND clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0004_
+ _0083_ Signal_Generator_1_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1162_ VGND VPWR VGND VPWR _0543_ _0531_ _0542_ _0544_ _0539_ sky130_fd_sc_hd__a2bb2o_1
X_1231_ VPWR VGND VGND VPWR _0595_ Dead_Time_Generator_inst_1.dt\[2\] _0596_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0601_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1093_ VPWR VGND VPWR VGND _0109_ _0499_ sky130_fd_sc_hd__inv_2
X_0877_ VPWR VGND _0054_ _0348_ Signal_Generator_2_90phase_inst.direction Signal_Generator_2_90phase_inst.count\[4\]
+ _0364_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0946_ VGND VPWR VGND VPWR _0414_ _0415_ _0410_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0731_ VPWR VGND VPWR VGND _0255_ _0241_ _0252_ _0003_ Signal_Generator_1_0phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0800_ VPWR VGND VGND VPWR _0304_ _0307_ _0020_ sky130_fd_sc_hd__nor2_1
X_0662_ VGND VPWR _0149_ _0205_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1214_ VGND VPWR _0588_ _0549_ _0545_ _0587_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1145_ VGND VPWR VGND VPWR Shift_Register_Inst.data_out\[13\] _0527_ net3 sky130_fd_sc_hd__or2b_1
X_1076_ VPWR VGND VPWR VGND _0094_ _0497_ sky130_fd_sc_hd__inv_2
X_0929_ VPWR VGND VGND VPWR _0404_ Signal_Generator_2_270phase_inst.count\[4\] _0390_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold46 net71 Signal_Generator_2_90phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net49 _0023_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net60 Signal_Generator_1_0phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 VPWR VGND VPWR VGND net38 Dead_Time_Generator_inst_1.dt\[3\] sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_7_Left_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0714_ VGND VPWR _0243_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ _0242_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0645_ VGND VPWR _0192_ _0194_ _0155_ _0188_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_1059_ VPWR VGND VPWR VGND _0078_ _0445_ sky130_fd_sc_hd__inv_2
X_1128_ VGND VPWR VPWR VGND _0510_ _0507_ _0502_ _0501_ _0508_ _0509_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput25 VPWR VGND VGND VPWR net25 SIGNAL_OUTPUT sky130_fd_sc_hd__buf_8
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0893_ VPWR VGND VPWR VGND _0376_ _0367_ _0374_ _0037_ net66 sky130_fd_sc_hd__a22o_1
X_0962_ VGND VPWR net17 _0425_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1161_ VPWR VGND VPWR VGND _0543_ net42 sky130_fd_sc_hd__inv_2
X_1230_ VPWR VGND VPWR VGND _0596_ Dead_Time_Generator_inst_1.dt\[2\] _0600_ _0597_
+ _0598_ _0599_ sky130_fd_sc_hd__a221o_1
X_1092_ VPWR VGND VPWR VGND _0108_ _0499_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ _0364_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0344_ Signal_Generator_2_90phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_42_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0945_ VGND VPWR VPWR VGND _0414_ net4 Shift_Register_Inst.data_out\[13\] _0413_
+ sky130_fd_sc_hd__mux2_1
X_1359_ Dead_Time_Generator_inst_2.count_dt\[2\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ _0166_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ VPWR VGND VPWR VGND _0254_ _0253_ _0244_ _0255_ sky130_fd_sc_hd__a21o_1
X_0661_ VGND VPWR VPWR VGND _0205_ Dead_Time_Generator_inst_1.dt\[3\] _0204_ _0182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1213_ VPWR VGND VGND VPWR _0585_ _0586_ _0587_ sky130_fd_sc_hd__nor2_1
X_1075_ VPWR VGND VPWR VGND _0093_ _0497_ sky130_fd_sc_hd__inv_2
X_1144_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[0\] _0503_ _0526_
+ _0523_ _0524_ _0525_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_23_Left_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0928_ VGND VPWR VPWR VGND Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0400_ _0403_ sky130_fd_sc_hd__or3b_1
X_0859_ VPWR VGND VGND VPWR _0351_ _0350_ _0347_ sky130_fd_sc_hd__or2_1
Xhold36 net61 Signal_Generator_2_90phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net72 Shift_Register_Inst.shift_state\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net50 Dead_Time_Generator_inst_1.count_dt\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net39 _0577_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0713_ VPWR VGND _0242_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
X_0644_ VPWR VGND VGND VPWR _0194_ _0191_ _0193_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1127_ VGND VPWR VGND VPWR Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[2\]
+ Shift_Register_Inst.data_out\[5\] Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[2\]
+ _0212_ _0509_ sky130_fd_sc_hd__mux4_1
X_1058_ VGND VPWR _0157_ _0496_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xoutput15 VGND VPWR net15 NMOS1_PS1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0961_ VPWR VGND _0425_ _0421_ _0416_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0892_ VPWR VGND VGND VPWR _0376_ _0370_ _0375_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1091_ VPWR VGND VPWR VGND _0107_ _0499_ sky130_fd_sc_hd__inv_2
X_1160_ VPWR VGND VPWR VGND _0540_ _0541_ _0539_ _0542_ sky130_fd_sc_hd__or3_1
X_0944_ VPWR VGND VPWR VGND _0413_ Dead_Time_Generator_inst_3.go sky130_fd_sc_hd__inv_2
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ VGND VPWR VPWR VGND _0053_ _0362_ _0361_ net77 _0346_ _0363_ sky130_fd_sc_hd__a32o_1
X_1358_ Dead_Time_Generator_inst_2.count_dt\[1\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ _0165_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1289_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0152_ _0073_ Shift_Register_Inst.shift_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0660_ VPWR VGND VGND VPWR _0204_ _0185_ _0191_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1212_ VPWR VGND VPWR VGND _0579_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_2.count_dt\[2\]
+ _0586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1074_ VPWR VGND VPWR VGND _0092_ _0497_ sky130_fd_sc_hd__inv_2
X_1143_ VGND VPWR _0525_ _0212_ _0208_ Signal_Generator_1_270phase_inst.count\[0\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_0927_ VPWR VGND VPWR VGND _0402_ _0388_ _0399_ _0045_ Signal_Generator_2_270phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ VPWR VGND VGND VPWR Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ _0350_ sky130_fd_sc_hd__nor2_1
X_0789_ VPWR VGND VGND VPWR _0299_ Signal_Generator_1_180phase_inst.count\[4\] _0285_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_15_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold26 net51 _0161_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 net73 _0198_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net40 _0582_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 net62 Dead_Time_Generator_inst_3.count_dt\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0712_ VGND VPWR VPWR VGND _0241_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0239_ _0240_ sky130_fd_sc_hd__o31a_2
X_0643_ VPWR VGND VGND VPWR _0188_ _0193_ Shift_Register_Inst.shift_state\[2\] sky130_fd_sc_hd__nand2_1
X_1126_ VGND VPWR VGND VPWR Shift_Register_Inst.data_out\[13\] _0508_ net5 sky130_fd_sc_hd__or2b_1
X_1057_ VGND VPWR _0496_ _0492_ _0456_ _0495_ VPWR VGND sky130_fd_sc_hd__and3_1
Xoutput16 VGND VPWR net16 NMOS1_PS2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1109_ VPWR VGND VPWR VGND _0124_ _0500_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0960_ VGND VPWR net22 _0424_ VPWR VGND sky130_fd_sc_hd__buf_1
X_0891_ VGND VPWR VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0375_ _0368_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1374_ Dead_Time_Generator_inst_3.go clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0181_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1090_ VPWR VGND VPWR VGND _0106_ _0499_ sky130_fd_sc_hd__inv_2
X_0874_ VGND VPWR _0344_ _0363_ Signal_Generator_2_90phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0943_ VGND VPWR net16 _0412_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0151_ _0072_ Dead_Time_Generator_inst_1.dt\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_1357_ Dead_Time_Generator_inst_2.count_dt\[0\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ _0164_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1142_ VPWR VGND VPWR VGND _0524_ Shift_Register_Inst.data_out\[6\] sky130_fd_sc_hd__inv_2
X_1211_ VGND VPWR _0585_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_2.count_dt\[2\]
+ _0579_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1073_ VPWR VGND VPWR VGND _0091_ _0497_ sky130_fd_sc_hd__inv_2
X_0926_ VPWR VGND VPWR VGND _0401_ _0400_ _0391_ _0402_ sky130_fd_sc_hd__a21o_1
X_0857_ VPWR VGND VPWR VGND _0049_ net61 sky130_fd_sc_hd__inv_2
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold38 net63 Signal_Generator_1_90phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ VGND VPWR VPWR VGND Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0295_ _0298_ sky130_fd_sc_hd__or3b_1
Xhold16 net41 Shift_Register_Inst.data_out\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 net52 Dead_Time_Generator_inst_1.count_dt\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net74 Signal_Generator_1_180phase_inst.direction VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ VPWR VGND VPWR VGND _0240_ Signal_Generator_1_0phase_inst.direction sky130_fd_sc_hd__inv_2
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR net26 clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
X_0642_ VPWR VGND VGND VPWR _0189_ _0191_ _0192_ sky130_fd_sc_hd__nor2_1
X_1125_ VPWR VGND VPWR VGND _0504_ _0507_ _0506_ Signal_Generator_1_180phase_inst.count\[3\]
+ _0503_ _0505_ sky130_fd_sc_hd__a2111o_1
X_1056_ VPWR VGND VPWR VGND _0480_ _0494_ _0468_ _0495_ sky130_fd_sc_hd__or3_1
X_0909_ VPWR VGND _0389_ Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[0\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_11_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput17 VGND VPWR net17 NMOS2_PS1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1108_ VPWR VGND VPWR VGND _0123_ _0500_ sky130_fd_sc_hd__inv_2
X_1039_ VGND VPWR _0478_ _0470_ net12 _0471_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_16_275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ VGND VPWR VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0374_ _0371_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1373_ Dead_Time_Generator_inst_4.count_dt\[4\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0180_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0873_ VPWR VGND VGND VPWR _0362_ Signal_Generator_2_90phase_inst.count\[4\] _0348_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_27_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0942_ VPWR VGND _0412_ _0411_ _0410_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_2_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1287_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0150_ _0071_ Dead_Time_Generator_inst_1.dt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_1356_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0163_ _0134_ Dead_Time_Generator_inst_1.dt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1141_ VGND VPWR VGND VPWR Signal_Generator_1_90phase_inst.count\[0\] _0523_ _0208_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ VPWR VGND VPWR VGND _0090_ _0497_ sky130_fd_sc_hd__inv_2
X_1210_ VGND VPWR _0165_ _0584_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0856_ VPWR VGND VGND VPWR _0346_ _0349_ _0055_ sky130_fd_sc_hd__nor2_1
X_0925_ VPWR VGND _0401_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_11_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0787_ VPWR VGND VPWR VGND _0297_ _0283_ _0294_ _0010_ net70 sky130_fd_sc_hd__a22o_1
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold28 net53 Dead_Time_Generator_inst_4.count_dt\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 net42 _0540_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net64 Dead_Time_Generator_inst_1.dt\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[1\] _0122_ _0036_
+ net29 sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0710_ VPWR VGND VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[0\]
+ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[3\]
+ _0239_ sky130_fd_sc_hd__or4_2
X_0641_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[1\] _0191_ _0190_ _0183_
+ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_27_Left_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1055_ VGND VPWR VPWR VGND _0493_ _0489_ _0486_ _0494_ sky130_fd_sc_hd__or3b_1
X_1124_ VPWR VGND VGND VPWR net44 _0212_ _0506_ sky130_fd_sc_hd__nor2_1
Xoutput18 VGND VPWR net18 NMOS2_PS2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0908_ _0388_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0386_ _0387_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_0839_ VPWR VGND VGND VPWR _0323_ _0336_ _0335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ VPWR VGND VPWR VGND _0122_ _0500_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1038_ VPWR VGND VGND VPWR _0472_ _0476_ _0477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1372_ Dead_Time_Generator_inst_4.count_dt\[3\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0179_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ VGND VPWR VPWR VGND _0411_ net5 Shift_Register_Inst.data_out\[13\] Dead_Time_Generator_inst_4.go
+ sky130_fd_sc_hd__mux2_1
X_0872_ VGND VPWR VPWR VGND Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0358_ _0361_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1355_ Dead_Time_Generator_inst_1.count_dt\[4\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0162_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1286_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0149_ _0070_ Dead_Time_Generator_inst_1.dt\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_41_Left_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1071_ VPWR VGND VPWR VGND _0089_ _0497_ sky130_fd_sc_hd__inv_2
X_1140_ VPWR VGND VGND VPWR _0000_ _0522_ _0506_ sky130_fd_sc_hd__nand2_1
X_0924_ VPWR VGND VPWR VGND _0400_ _0390_ sky130_fd_sc_hd__inv_2
X_0855_ VGND VPWR _0349_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.count\[5\]
+ _0348_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0786_ VPWR VGND VPWR VGND _0296_ _0295_ _0286_ _0297_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1338_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[0\] _0121_ _0035_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold18 net43 _0159_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net54 Signal_Generator_2_0phase_inst.count\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ VGND VPWR _0629_ _0495_ _0492_ _0628_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_29_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0640_ VPWR VGND VPWR VGND _0190_ Shift_Register_Inst.shift_state\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_20_185 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1054_ VPWR VGND _0493_ _0487_ _0488_ VPWR VGND sky130_fd_sc_hd__and2_1
X_1123_ VGND VPWR _0505_ Shift_Register_Inst.data_out\[6\] Shift_Register_Inst.data_out\[5\]
+ Signal_Generator_1_270phase_inst.count\[3\] VPWR VGND sky130_fd_sc_hd__and3_1
X_0907_ VPWR VGND VPWR VGND _0387_ Signal_Generator_2_270phase_inst.direction sky130_fd_sc_hd__inv_2
XFILLER_0_28_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput19 VGND VPWR net19 NMOS_PS3 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0838_ VPWR VGND Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] _0335_ Signal_Generator_2_0phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0769_ VPWR VGND _0284_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_44_Left_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1106_ VPWR VGND VPWR VGND _0121_ _0500_ sky130_fd_sc_hd__inv_2
X_1037_ VPWR VGND VPWR VGND _0475_ _0474_ net11 _0476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ Dead_Time_Generator_inst_4.count_dt\[2\] clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ _0178_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0940_ VPWR VGND VGND VPWR Shift_Register_Inst.data_out\[17\] Shift_Register_Inst.data_out\[16\]
+ _0410_ Shift_Register_Inst.data_out\[15\] sky130_fd_sc_hd__nor3b_1
X_0871_ VPWR VGND VPWR VGND _0360_ _0346_ _0357_ _0052_ net71 sky130_fd_sc_hd__a22o_1
X_1354_ Dead_Time_Generator_inst_1.count_dt\[3\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ net51 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1285_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0148_ _0069_ Dead_Time_Generator_inst_1.dt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_60 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ VPWR VGND VPWR VGND _0088_ _0497_ sky130_fd_sc_hd__inv_2
X_0923_ VPWR VGND VGND VPWR _0386_ _0399_ _0398_ sky130_fd_sc_hd__nand2_1
X_0854_ VGND VPWR _0348_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ _0347_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0785_ VPWR VGND _0296_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_23_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1337_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.direction _0120_ _0041_
+ net29 sky130_fd_sc_hd__dfstp_2
X_1268_ VPWR VGND VPWR VGND _0622_ Dead_Time_Generator_inst_4.count_dt\[3\] Dead_Time_Generator_inst_4.count_dt\[4\]
+ _0628_ sky130_fd_sc_hd__a21o_1
Xhold19 net44 Shift_Register_Inst.data_out\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1199_ VPWR VGND VGND VPWR _0569_ Dead_Time_Generator_inst_1.dt\[2\] _0570_ net38
+ _0575_ sky130_fd_sc_hd__o22a_1
X_1122_ Shift_Register_Inst.data_out\[6\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0504_ Shift_Register_Inst.data_out\[5\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_1053_ VPWR VGND VGND VPWR _0465_ _0466_ _0492_ _0491_ _0468_ sky130_fd_sc_hd__o22ai_2
X_0906_ VPWR VGND VPWR VGND Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[2\]
+ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[0\]
+ _0386_ sky130_fd_sc_hd__or4_2
X_0837_ VPWR VGND VPWR VGND _0334_ _0325_ _0332_ _0030_ Signal_Generator_2_0phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0768_ VGND VPWR VPWR VGND _0283_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0281_ _0282_ sky130_fd_sc_hd__o31a_2
X_0699_ VGND VPWR VPWR VGND _0232_ Shift_Register_Inst.data_out\[14\] _0231_ net1
+ sky130_fd_sc_hd__mux2_1
X_1105_ VPWR VGND VPWR VGND _0120_ _0500_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1036_ VPWR VGND VGND VPWR Signal_Generator_2_0phase_inst.count\[2\] _0475_ _0458_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ VPWR VGND VGND VPWR _0217_ _0458_ _0215_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ Dead_Time_Generator_inst_4.count_dt\[1\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0177_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ VPWR VGND VPWR VGND _0359_ _0358_ _0349_ _0360_ sky130_fd_sc_hd__a21o_1
Xclkbuf_3_2__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_1284_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0147_ _0068_ Shift_Register_Inst.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_1353_ Dead_Time_Generator_inst_1.count_dt\[2\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ _0160_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0999_ VPWR VGND VPWR VGND _0071_ _0444_ sky130_fd_sc_hd__inv_2
X_0922_ VPWR VGND Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] _0398_ Signal_Generator_2_270phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0853_ VPWR VGND _0347_ Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[0\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
X_0784_ VPWR VGND VPWR VGND _0295_ _0285_ sky130_fd_sc_hd__inv_2
X_1336_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0054_
+ _0119_ Signal_Generator_2_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1267_ VGND VPWR _0179_ _0627_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xinput1 VPWR VGND net1 Data_SR VPWR VGND sky130_fd_sc_hd__buf_2
X_1198_ VPWR VGND VPWR VGND _0570_ Dead_Time_Generator_inst_1.dt\[2\] _0574_ _0571_
+ _0572_ _0573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1052_ VPWR VGND VGND VPWR _0490_ _0478_ _0477_ _0480_ _0491_ sky130_fd_sc_hd__o22a_1
X_1121_ _0503_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0905_ VPWR VGND _0040_ _0369_ Signal_Generator_2_180phase_inst.direction Signal_Generator_2_180phase_inst.count\[4\]
+ _0385_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0767_ VPWR VGND VPWR VGND _0282_ Signal_Generator_1_180phase_inst.direction sky130_fd_sc_hd__inv_2
X_0836_ VPWR VGND VGND VPWR _0334_ _0328_ _0333_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0698_ VPWR VGND VGND VPWR _0231_ _0228_ _0201_ sky130_fd_sc_hd__or2_1
X_1319_ VGND VPWR VPWR VGND clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0016_
+ _0102_ Signal_Generator_1_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1104_ VPWR VGND VPWR VGND _0119_ _0500_ sky130_fd_sc_hd__inv_2
X_1035_ VGND VPWR VGND VPWR _0459_ Signal_Generator_2_180phase_inst.count\[2\] _0460_
+ Signal_Generator_2_90phase_inst.count\[2\] _0474_ _0473_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_3_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ VGND VPWR VPWR VGND _0018_ _0320_ _0319_ Signal_Generator_1_270phase_inst.direction
+ _0304_ _0321_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1018_ VPWR VGND _0457_ _0217_ _0215_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_19 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1283_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0146_ _0067_ Shift_Register_Inst.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_1352_ Dead_Time_Generator_inst_1.count_dt\[1\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ net43 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0998_ VPWR VGND VPWR VGND _0070_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0921_ VPWR VGND VPWR VGND _0397_ _0388_ _0395_ _0044_ Signal_Generator_2_270phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0852_ VGND VPWR VPWR VGND _0346_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0344_ _0345_ sky130_fd_sc_hd__o31a_2
X_0783_ VPWR VGND VGND VPWR _0281_ _0294_ _0293_ sky130_fd_sc_hd__nand2_1
X_1335_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[4\] _0118_ _0053_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
X_1266_ VGND VPWR _0627_ _0594_ _0593_ _0626_ VPWR VGND sky130_fd_sc_hd__and3_1
Xinput2 VGND VPWR net2 net37 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1197_ _0573_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_14_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1051_ VPWR VGND VGND VPWR _0486_ _0489_ _0490_ sky130_fd_sc_hd__nor2_1
X_1120_ VPWR VGND VPWR VGND _0212_ Signal_Generator_1_0phase_inst.count\[3\] _0208_
+ _0502_ sky130_fd_sc_hd__or3_1
X_0904_ _0385_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0365_ Signal_Generator_2_180phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0766_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[0\]
+ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[3\]
+ _0281_ sky130_fd_sc_hd__or4_2
X_0697_ VGND VPWR _0139_ _0230_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0835_ VGND VPWR VPWR VGND Signal_Generator_2_0phase_inst.count\[2\] _0333_ _0326_
+ sky130_fd_sc_hd__xor2_1
X_1318_ VGND VPWR VPWR VGND clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0015_
+ _0101_ Signal_Generator_1_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1249_ VPWR VGND VGND VPWR _0577_ _0614_ _0578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1103_ VPWR VGND VPWR VGND _0118_ _0500_ sky130_fd_sc_hd__inv_2
X_1034_ VGND VPWR _0473_ _0217_ _0215_ Signal_Generator_2_270phase_inst.count\[2\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_17_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0749_ VPWR VGND VPWR VGND _0268_ _0262_ _0267_ _0022_ Signal_Generator_1_90phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0818_ VGND VPWR _0302_ _0321_ Signal_Generator_1_270phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_32_Left_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1017_ VPWR VGND VGND VPWR _0454_ _0456_ _0455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1351_ Dead_Time_Generator_inst_1.count_dt\[0\] clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ net33 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1282_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0145_ _0066_ Shift_Register_Inst.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ VPWR VGND VPWR VGND _0069_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0920_ VPWR VGND VGND VPWR _0397_ _0391_ _0396_ sky130_fd_sc_hd__or2_1
X_0851_ VPWR VGND VPWR VGND _0345_ Signal_Generator_2_90phase_inst.direction sky130_fd_sc_hd__inv_2
X_0782_ VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] _0293_ Signal_Generator_1_180phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_1334_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[3\] _0117_ _0052_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1265_ VGND VPWR _0622_ _0626_ _0446_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1196_ _0572_ Dead_Time_Generator_inst_2.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xinput3 VGND VPWR net3 d1[0] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1050_ VGND VPWR VPWR VGND _0489_ net10 _0485_ _0488_ _0487_ sky130_fd_sc_hd__o2bb2a_1
X_0903_ VGND VPWR VPWR VGND _0039_ _0383_ _0382_ Signal_Generator_2_180phase_inst.direction
+ _0367_ _0384_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0834_ VGND VPWR VPWR VGND Signal_Generator_2_0phase_inst.count\[2\] _0332_ _0329_
+ sky130_fd_sc_hd__xor2_1
X_0765_ VPWR VGND _0026_ _0264_ Signal_Generator_1_90phase_inst.direction Signal_Generator_1_90phase_inst.count\[4\]
+ _0280_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0696_ VGND VPWR VPWR VGND _0230_ Shift_Register_Inst.data_out\[13\] _0229_ net1
+ sky130_fd_sc_hd__mux2_1
X_1317_ VGND VPWR VPWR VGND clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0014_
+ _0100_ Signal_Generator_1_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1248_ VGND VPWR VPWR VGND _0174_ _0593_ _0594_ net59 _0612_ sky130_fd_sc_hd__o2bb2a_1
X_1179_ VPWR VGND _0561_ net31 _0558_ VPWR VGND sky130_fd_sc_hd__and2_1
X_1102_ VPWR VGND VPWR VGND _0117_ _0500_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ VPWR VGND VPWR VGND _0471_ _0470_ net12 _0472_ sky130_fd_sc_hd__a21oi_1
X_0817_ VPWR VGND VGND VPWR _0320_ Signal_Generator_1_270phase_inst.count\[4\] _0306_
+ sky130_fd_sc_hd__or2_1
X_0748_ VGND VPWR VGND VPWR _0265_ _0268_ _0267_ sky130_fd_sc_hd__or2b_1
X_0679_ VPWR VGND VPWR VGND _0188_ _0184_ Shift_Register_Inst.shift_state\[2\] _0183_
+ _0218_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ VGND VPWR VGND VPWR net30 _0455_ Dead_Time_Generator_inst_4.count_dt\[4\]
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_62 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1350_ VPWR VGND VPWR VGND Signal_Generator_2_270phase_inst.count\[5\] _0133_ _0047_
+ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1281_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0144_ _0065_ Shift_Register_Inst.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_0996_ VPWR VGND VPWR VGND _0068_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[2\]
+ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[0\]
+ _0344_ sky130_fd_sc_hd__or4_2
X_0781_ VPWR VGND VPWR VGND _0292_ _0283_ _0290_ _0009_ net70 sky130_fd_sc_hd__a22o_1
X_1333_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0116_ _0051_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
X_1264_ VGND VPWR _0178_ _0625_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xinput4 VGND VPWR net4 d1[1] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1195_ VGND VPWR VGND VPWR Dead_Time_Generator_inst_1.dt\[1\] _0571_ Dead_Time_Generator_inst_2.count_dt\[1\]
+ sky130_fd_sc_hd__or2b_1
X_0979_ VGND VPWR VGND VPWR _0440_ _0434_ net25 _0427_ sky130_fd_sc_hd__a21bo_4
X_0902_ VGND VPWR _0365_ _0384_ Signal_Generator_2_180phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0833_ VPWR VGND VPWR VGND _0331_ _0325_ _0330_ _0029_ Signal_Generator_2_0phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0764_ _0280_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0260_ Signal_Generator_1_90phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_0695_ VPWR VGND VGND VPWR _0229_ _0228_ _0209_ sky130_fd_sc_hd__or2_1
X_1247_ VPWR VGND VPWR VGND _0173_ _0613_ _0612_ _0593_ _0594_ sky130_fd_sc_hd__a211oi_1
X_1178_ VGND VPWR _0560_ _0558_ Dead_Time_Generator_inst_1.count_dt\[0\] net31 VPWR
+ VGND sky130_fd_sc_hd__and3_1
X_1316_ VGND VPWR VPWR VGND clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0020_
+ _0099_ Signal_Generator_1_270phase_inst.direction sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1101_ VPWR VGND VPWR VGND _0116_ _0500_ sky130_fd_sc_hd__inv_2
X_1032_ VPWR VGND VGND VPWR Signal_Generator_2_0phase_inst.count\[3\] _0471_ _0458_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0747_ VPWR VGND VGND VPWR _0267_ _0266_ _0263_ sky130_fd_sc_hd__or2_1
X_0816_ VGND VPWR VPWR VGND Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0316_ _0319_ sky130_fd_sc_hd__or3b_1
X_0678_ VPWR VGND _0217_ Shift_Register_Inst.data_out\[8\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1015_ VPWR VGND VPWR VGND _0446_ net38 _0454_ _0451_ _0452_ _0453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1280_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0143_ _0064_ Shift_Register_Inst.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_0995_ VPWR VGND VPWR VGND _0067_ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ VPWR VGND VGND VPWR _0292_ _0286_ _0291_ sky130_fd_sc_hd__or2_1
X_1332_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[1\] _0115_ _0050_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1263_ VGND VPWR _0625_ _0594_ _0593_ _0624_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1194_ VPWR VGND VPWR VGND _0570_ Dead_Time_Generator_inst_2.count_dt\[2\] sky130_fd_sc_hd__inv_2
Xinput5 VGND VPWR net5 d1[2] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ VGND VPWR VGND VPWR _0439_ Shift_Register_Inst.data_out\[9\] _0436_ _0427_
+ Shift_Register_Inst.data_out\[11\] _0440_ sky130_fd_sc_hd__o32a_2
XFILLER_0_9_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0901_ VPWR VGND VGND VPWR _0383_ Signal_Generator_2_180phase_inst.count\[4\] _0369_
+ sky130_fd_sc_hd__or2_1
X_0763_ VGND VPWR VPWR VGND _0025_ _0278_ _0277_ Signal_Generator_1_90phase_inst.direction
+ _0262_ _0279_ sky130_fd_sc_hd__a32o_1
X_0832_ VGND VPWR VGND VPWR _0328_ _0331_ _0330_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1315_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[5\] _0098_ _0012_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_0694_ VPWR VGND VGND VPWR Shift_Register_Inst.shift_state\[3\] _0228_ Shift_Register_Inst.shift_state\[2\]
+ sky130_fd_sc_hd__nand2_1
X_1177_ VGND VPWR VGND VPWR net30 _0559_ Dead_Time_Generator_inst_1.count_dt\[4\]
+ sky130_fd_sc_hd__or2b_1
X_1246_ VPWR VGND VGND VPWR _0596_ _0608_ _0595_ _0613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ VGND VPWR VGND VPWR _0459_ Signal_Generator_2_180phase_inst.count\[3\] _0460_
+ Signal_Generator_2_90phase_inst.count\[3\] _0470_ _0469_ sky130_fd_sc_hd__a221oi_2
X_1100_ VPWR VGND _0500_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_33_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0746_ VPWR VGND VGND VPWR net47 Signal_Generator_1_90phase_inst.count\[0\] _0266_
+ sky130_fd_sc_hd__nor2_1
X_0815_ VPWR VGND VPWR VGND _0318_ _0304_ _0315_ _0017_ net80 sky130_fd_sc_hd__a22o_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0677_ VGND VPWR _0145_ _0216_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1229_ _0599_ Dead_Time_Generator_inst_3.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_0_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0453_ Dead_Time_Generator_inst_4.count_dt\[4\] Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_8_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ VPWR VGND _0254_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_45_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ VPWR VGND VPWR VGND _0066_ _0444_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Left_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1331_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.count\[0\] _0114_ _0049_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1262_ VPWR VGND VGND VPWR _0622_ _0623_ _0624_ sky130_fd_sc_hd__nor2_1
X_1193_ VPWR VGND VPWR VGND _0569_ Dead_Time_Generator_inst_2.count_dt\[3\] sky130_fd_sc_hd__inv_2
Xinput6 VGND VPWR net6 d1[3] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ VPWR VGND VGND VPWR _0439_ _0438_ Shift_Register_Inst.data_out\[10\] sky130_fd_sc_hd__nand2_2
XFILLER_0_9_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0900_ VGND VPWR VPWR VGND Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0379_ _0382_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0762_ VGND VPWR _0260_ _0279_ Signal_Generator_1_90phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_0693_ VGND VPWR _0140_ _0227_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0831_ VPWR VGND VGND VPWR _0330_ _0329_ _0326_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1314_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[4\] _0097_ _0011_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
Xclkbuf_0_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR Dead_Time_Generator_inst_1.clk
+ clknet_0_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_1176_ VPWR VGND VPWR VGND _0550_ net67 _0558_ _0555_ _0556_ _0557_ sky130_fd_sc_hd__a221o_1
X_1245_ _0612_ Dead_Time_Generator_inst_3.count_dt\[1\] Dead_Time_Generator_inst_3.count_dt\[3\]
+ Dead_Time_Generator_inst_3.count_dt\[2\] _0605_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_6_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1030_ VGND VPWR _0469_ _0217_ _0215_ Signal_Generator_2_270phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_0814_ VPWR VGND VPWR VGND _0317_ _0316_ _0307_ _0318_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_26_Left_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0745_ VPWR VGND VPWR VGND _0021_ net63 sky130_fd_sc_hd__inv_2
X_0676_ VGND VPWR VPWR VGND _0216_ _0215_ _0194_ _0182_ sky130_fd_sc_hd__mux2_1
X_1228_ _0598_ Dead_Time_Generator_inst_3.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_1159_ VPWR VGND VGND VPWR _0532_ _0533_ _0541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1013_ VPWR VGND VGND VPWR _0446_ Dead_Time_Generator_inst_1.dt\[2\] _0447_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0452_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0728_ VPWR VGND VPWR VGND _0253_ _0243_ sky130_fd_sc_hd__inv_2
X_0659_ VGND VPWR _0150_ _0203_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Left_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0993_ VPWR VGND _0444_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_41_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ VPWR VGND VPWR VGND Signal_Generator_2_90phase_inst.direction _0113_ _0055_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1261_ VPWR VGND VPWR VGND _0616_ net53 Dead_Time_Generator_inst_4.count_dt\[2\]
+ _0623_ sky130_fd_sc_hd__a21oi_1
Xinput7 VGND VPWR net7 d1[4] VPWR VGND sky130_fd_sc_hd__buf_1
X_1192_ VPWR VGND VPWR VGND _0134_ _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0976_ VGND VPWR VGND VPWR _0438_ _0437_ _0427_ Shift_Register_Inst.data_out\[11\]
+ net23 sky130_fd_sc_hd__a31o_4
XPHY_EDGE_ROW_40_Left_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ VPWR VGND VGND VPWR Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ _0329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0761_ VPWR VGND VGND VPWR _0278_ Signal_Generator_1_90phase_inst.count\[4\] _0264_
+ sky130_fd_sc_hd__or2_1
X_0692_ VGND VPWR VPWR VGND _0227_ Shift_Register_Inst.data_out\[12\] _0226_ net1
+ sky130_fd_sc_hd__mux2_1
X_1313_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[3\] _0096_ _0010_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1244_ VPWR VGND VPWR VGND _0594_ _0593_ _0611_ _0172_ sky130_fd_sc_hd__a21oi_1
X_1175_ _0557_ Dead_Time_Generator_inst_1.count_dt\[4\] net30 VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0959_ VPWR VGND VGND VPWR _0424_ _0414_ _0423_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xinput10 VGND VPWR net10 d2[1] VPWR VGND sky130_fd_sc_hd__buf_1
X_0813_ VPWR VGND _0317_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0675_ VGND VPWR Shift_Register_Inst.data_out\[7\] _0215_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_0744_ VPWR VGND VGND VPWR _0262_ net35 _0027_ sky130_fd_sc_hd__nor2_1
X_1158_ VPWR VGND VGND VPWR _0534_ _0538_ _0540_ sky130_fd_sc_hd__nor2_1
X_1227_ VGND VPWR VGND VPWR Dead_Time_Generator_inst_1.dt\[1\] _0597_ Dead_Time_Generator_inst_3.count_dt\[1\]
+ sky130_fd_sc_hd__or2b_1
X_1089_ VPWR VGND _0499_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_30_222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1012_ VPWR VGND VPWR VGND _0447_ Dead_Time_Generator_inst_1.dt\[2\] _0451_ _0448_
+ _0449_ _0450_ sky130_fd_sc_hd__a221o_1
X_0727_ VPWR VGND VGND VPWR _0239_ _0252_ _0251_ sky130_fd_sc_hd__nand2_1
X_0658_ VGND VPWR VPWR VGND _0203_ Dead_Time_Generator_inst_1.dt\[2\] _0202_ _0182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_185 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ VPWR VGND VPWR VGND _0065_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ VGND VPWR _0622_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_4.count_dt\[2\]
+ _0616_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_36_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 VGND VPWR net8 d1[5] VPWR VGND sky130_fd_sc_hd__buf_1
X_1191_ VGND VPWR VPWR VGND _0162_ _0545_ _0549_ net55 _0567_ sky130_fd_sc_hd__o2bb2a_1
X_0975_ VGND VPWR VGND VPWR _0437_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ Shift_Register_Inst.data_out\[12\] Shift_Register_Inst.data_out\[11\] sky130_fd_sc_hd__and3b_2
Xclkbuf_3_4__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR net28 clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0760_ VGND VPWR VPWR VGND Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0274_ _0277_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0691_ VPWR VGND VPWR VGND _0188_ _0184_ _0189_ _0183_ _0226_ sky130_fd_sc_hd__or4_1
X_1312_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0095_ _0009_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
X_1174_ VPWR VGND VGND VPWR _0550_ Dead_Time_Generator_inst_1.dt\[2\] _0551_ Dead_Time_Generator_inst_1.dt\[3\]
+ _0556_ sky130_fd_sc_hd__o22a_1
X_1243_ VGND VPWR _0608_ _0611_ _0596_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0889_ VPWR VGND VPWR VGND _0373_ _0367_ _0372_ _0036_ Signal_Generator_2_180phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ VPWR VGND VGND VPWR _0423_ Shift_Register_Inst.data_out\[17\] Shift_Register_Inst.data_out\[15\]
+ Shift_Register_Inst.data_out\[16\] sky130_fd_sc_hd__nand3b_1
XFILLER_0_33_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 VGND VPWR net11 d2[2] VPWR VGND sky130_fd_sc_hd__buf_1
X_0743_ VGND VPWR _0265_ Signal_Generator_1_90phase_inst.count\[4\] net34 _0264_ VPWR
+ VGND sky130_fd_sc_hd__and3_1
X_0812_ VPWR VGND VPWR VGND _0316_ _0306_ sky130_fd_sc_hd__inv_2
X_0674_ VGND VPWR _0146_ _0214_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1157_ VPWR VGND VPWR VGND _0534_ _0532_ _0533_ _0539_ _0538_ sky130_fd_sc_hd__a22o_1
X_1226_ VPWR VGND VPWR VGND _0596_ net75 sky130_fd_sc_hd__inv_2
X_1088_ VPWR VGND VPWR VGND _0105_ _0498_ sky130_fd_sc_hd__inv_2
X_1011_ _0450_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0726_ VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] _0251_ Signal_Generator_1_0phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0657_ VPWR VGND VGND VPWR _0202_ _0185_ _0201_ sky130_fd_sc_hd__or2_1
X_1209_ VGND VPWR _0584_ _0549_ _0545_ _0583_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ VGND VPWR _0135_ _0238_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ VPWR VGND VPWR VGND _0064_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ VPWR VGND VPWR VGND _0161_ _0568_ _0567_ _0545_ _0549_ sky130_fd_sc_hd__a211oi_1
Xinput9 VGND VPWR net9 d2[0] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0974_ VPWR VGND VPWR VGND _0430_ net24 _0435_ _0436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0690_ VGND VPWR _0141_ _0225_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1311_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[1\] _0094_ _0008_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
X_1242_ VPWR VGND VPWR VGND _0594_ _0593_ _0610_ _0171_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1173_ VPWR VGND VPWR VGND _0551_ Dead_Time_Generator_inst_1.dt\[2\] _0555_ _0552_
+ _0553_ _0554_ sky130_fd_sc_hd__a221o_1
X_0888_ VGND VPWR VGND VPWR _0370_ _0373_ _0372_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ VGND VPWR net15 _0422_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput12 VGND VPWR net12 d2[3] VPWR VGND sky130_fd_sc_hd__buf_1
X_0742_ VGND VPWR _0264_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0263_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0811_ VPWR VGND VGND VPWR _0302_ _0315_ _0314_ sky130_fd_sc_hd__nand2_1
X_0673_ VGND VPWR VPWR VGND _0214_ _0212_ _0213_ _0182_ sky130_fd_sc_hd__mux2_1
X_1225_ VPWR VGND VPWR VGND _0595_ net68 sky130_fd_sc_hd__inv_2
X_1156_ VGND VPWR VGND VPWR _0538_ _0506_ _0535_ Signal_Generator_1_0phase_inst.count\[5\]
+ _0537_ sky130_fd_sc_hd__a211o_1
X_1087_ VPWR VGND VPWR VGND _0104_ _0498_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1010_ _0449_ Dead_Time_Generator_inst_4.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0725_ VPWR VGND VPWR VGND _0250_ _0241_ _0248_ _0002_ net78 sky130_fd_sc_hd__a22o_1
X_0656_ VGND VPWR VPWR VGND Shift_Register_Inst.shift_state\[0\] Shift_Register_Inst.shift_state\[1\]
+ _0183_ _0201_ sky130_fd_sc_hd__or3b_1
X_1208_ VGND VPWR VPWR VGND Dead_Time_Generator_inst_2.count_dt\[1\] _0583_ _0579_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1139_ VPWR VGND VGND VPWR _0521_ _0519_ _0520_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0708_ VGND VPWR VPWR VGND _0238_ Shift_Register_Inst.data_out\[17\] _0237_ net1
+ sky130_fd_sc_hd__mux2_1
X_0639_ VPWR VGND VPWR VGND _0189_ Shift_Register_Inst.shift_state\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0990_ VPWR VGND VPWR VGND _0063_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0973_ VGND VPWR _0435_ _0428_ Shift_Register_Inst.data_out\[9\] net19 VPWR VGND
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Left_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1241_ VPWR VGND VGND VPWR _0608_ _0610_ _0609_ sky130_fd_sc_hd__nand2_1
X_1310_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.count\[0\] _0093_ _0007_
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0554_ Dead_Time_Generator_inst_1.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_42_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0956_ VPWR VGND _0422_ _0421_ _0411_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0887_ VPWR VGND VGND VPWR _0372_ _0371_ _0368_ sky130_fd_sc_hd__or2_1
Xinput13 VGND VPWR net13 d2[4] VPWR VGND sky130_fd_sc_hd__buf_1
X_0810_ VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] _0314_ Signal_Generator_1_270phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0741_ VPWR VGND _0263_ Signal_Generator_1_90phase_inst.count\[0\] net47 VPWR VGND
+ sky130_fd_sc_hd__and2_1
X_0672_ VPWR VGND VGND VPWR _0213_ _0193_ _0201_ sky130_fd_sc_hd__or2_1
X_1224_ VPWR VGND _0594_ _0495_ VPWR VGND sky130_fd_sc_hd__buf_2
X_1155_ VPWR VGND VPWR VGND _0503_ Signal_Generator_1_180phase_inst.count\[5\] _0536_
+ _0537_ sky130_fd_sc_hd__a21o_1
X_1086_ VPWR VGND VPWR VGND _0103_ _0498_ sky130_fd_sc_hd__inv_2
X_0939_ VPWR VGND VGND VPWR net24 Shift_Register_Inst.data_out\[16\] _0409_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_5_Left_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0724_ VPWR VGND VGND VPWR _0250_ _0244_ _0249_ sky130_fd_sc_hd__or2_1
X_0655_ VGND VPWR _0151_ _0200_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1207_ VGND VPWR _0164_ net40 VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1069_ VPWR VGND VPWR VGND _0087_ _0497_ sky130_fd_sc_hd__inv_2
X_1138_ VGND VPWR VGND VPWR Shift_Register_Inst.data_out\[13\] _0520_ net4 sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_31_Left_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ VPWR VGND VPWR VGND _0190_ _0185_ Shift_Register_Inst.shift_state\[1\] _0237_
+ _0183_ sky130_fd_sc_hd__or4b_1
X_0638_ VPWR VGND VPWR VGND _0188_ Shift_Register_Inst.shift_state\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ VGND VPWR VPWR VGND _0434_ _0433_ Shift_Register_Inst.data_out\[11\] _0429_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ _0553_ Dead_Time_Generator_inst_1.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_1240_ VPWR VGND VGND VPWR _0609_ Dead_Time_Generator_inst_3.count_dt\[1\] _0605_
+ sky130_fd_sc_hd__or2_1
X_0886_ VPWR VGND VGND VPWR net65 Signal_Generator_2_180phase_inst.count\[1\] _0371_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0955_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] _0421_
+ Shift_Register_Inst.data_out\[15\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ Dead_Time_Generator_inst_4.count_dt\[0\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0176_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xinput14 VGND VPWR net14 d2[5] VPWR VGND sky130_fd_sc_hd__buf_1
X_0740_ _0262_ net34 Signal_Generator_1_90phase_inst.count\[4\] _0260_ _0261_ VPWR
+ VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_3_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0671_ VPWR VGND _0212_ Shift_Register_Inst.data_out\[6\] VPWR VGND sky130_fd_sc_hd__buf_2
X_1223_ VPWR VGND _0593_ _0492_ VPWR VGND sky130_fd_sc_hd__buf_2
X_1154_ VGND VPWR _0536_ Shift_Register_Inst.data_out\[6\] Shift_Register_Inst.data_out\[5\]
+ Signal_Generator_1_270phase_inst.count\[5\] VPWR VGND sky130_fd_sc_hd__and3_1
X_1085_ VPWR VGND VPWR VGND _0102_ _0498_ sky130_fd_sc_hd__inv_2
X_0869_ VPWR VGND _0359_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0938_ VPWR VGND VPWR VGND _0409_ net7 sky130_fd_sc_hd__inv_2
XFILLER_0_3_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ VGND VPWR VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] _0249_ _0242_
+ sky130_fd_sc_hd__xor2_1
X_0654_ VGND VPWR VPWR VGND _0200_ Dead_Time_Generator_inst_1.dt\[1\] _0199_ _0182_
+ sky130_fd_sc_hd__mux2_1
X_1137_ VPWR VGND VGND VPWR _0519_ _0518_ _0517_ _0516_ _0515_ _0506_ sky130_fd_sc_hd__o41a_1
X_1206_ VGND VPWR _0582_ _0549_ _0545_ _0581_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1068_ VPWR VGND VPWR VGND _0086_ _0497_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0706_ VGND VPWR _0136_ _0236_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0637_ VGND VPWR Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ Shift_Register_Inst.shift_state\[2\] _0156_ _0183_ net76 VPWR VGND sky130_fd_sc_hd__a41o_1
Xclkbuf_3_5__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk
+ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0971_ VPWR VGND VPWR VGND net21 _0430_ _0433_ _0431_ net16 _0432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ VGND VPWR VGND VPWR Dead_Time_Generator_inst_1.dt\[1\] _0552_ Dead_Time_Generator_inst_1.count_dt\[1\]
+ sky130_fd_sc_hd__or2b_1
X_0885_ VPWR VGND VPWR VGND _0035_ net65 sky130_fd_sc_hd__inv_2
XFILLER_0_27_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ VGND VPWR net21 _0420_ VPWR VGND sky130_fd_sc_hd__buf_1
X_1299_ VGND VPWR VPWR VGND clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0003_
+ _0082_ Signal_Generator_1_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1368_ Dead_Time_Generator_inst_2.go clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0175_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0670_ VGND VPWR _0147_ _0211_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1153_ VGND VPWR _0535_ _0524_ _0208_ Signal_Generator_1_90phase_inst.count\[5\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_1222_ VPWR VGND VPWR VGND _0549_ _0545_ _0561_ _0169_ sky130_fd_sc_hd__a21oi_1
X_1084_ VPWR VGND VPWR VGND _0101_ _0498_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0868_ VPWR VGND VPWR VGND _0358_ _0348_ sky130_fd_sc_hd__inv_2
X_0799_ VGND VPWR _0307_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.count\[5\]
+ _0306_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0937_ VPWR VGND VPWR VGND net19 _0408_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0722_ VGND VPWR VPWR VGND Signal_Generator_1_0phase_inst.count\[2\] _0248_ _0245_
+ sky130_fd_sc_hd__xor2_1
X_0653_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[1\] _0185_ _0190_ _0183_
+ _0199_ sky130_fd_sc_hd__or4_1
X_1067_ VPWR VGND _0497_ _0441_ VPWR VGND sky130_fd_sc_hd__buf_4
X_1136_ VPWR VGND VPWR VGND _0212_ Signal_Generator_1_0phase_inst.count\[1\] _0208_
+ _0518_ sky130_fd_sc_hd__or3_1
X_1205_ VPWR VGND VGND VPWR _0579_ _0580_ _0581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0705_ VGND VPWR VPWR VGND _0236_ Shift_Register_Inst.data_out\[16\] _0235_ net1
+ sky130_fd_sc_hd__mux2_1
X_0636_ VGND VPWR _0163_ _0187_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1119_ VGND VPWR VGND VPWR Shift_Register_Inst.data_out\[13\] _0501_ net6 sky130_fd_sc_hd__or2b_1
XFILLER_0_28_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0970_ VGND VPWR _0432_ _0428_ Shift_Register_Inst.data_out\[9\] net18 VPWR VGND
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0884_ VPWR VGND VGND VPWR _0367_ _0370_ _0041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_255 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0953_ VGND VPWR VGND VPWR _0419_ _0420_ _0410_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ Dead_Time_Generator_inst_3.count_dt\[4\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0174_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1298_ VGND VPWR VPWR VGND clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0002_
+ _0081_ Signal_Generator_1_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_236 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1221_ VGND VPWR _0168_ _0592_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f_CLK_SR VGND VPWR VGND VPWR clknet_0_CLK_SR clknet_1_1__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
X_1152_ VGND VPWR VGND VPWR net41 _0534_ net8 sky130_fd_sc_hd__or2b_1
X_1083_ VPWR VGND VPWR VGND _0100_ _0498_ sky130_fd_sc_hd__inv_2
X_0936_ VPWR VGND _0408_ net8 Shift_Register_Inst.data_out\[16\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_23_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0867_ VPWR VGND VGND VPWR _0344_ _0357_ _0356_ sky130_fd_sc_hd__nand2_1
X_0798_ VGND VPWR _0306_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ _0305_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_15_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0721_ VPWR VGND VPWR VGND _0247_ _0241_ _0246_ _0001_ Signal_Generator_1_0phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0652_ VPWR VGND VGND VPWR _0197_ net73 _0152_ sky130_fd_sc_hd__nor2_1
X_1204_ VPWR VGND VPWR VGND _0578_ net39 Dead_Time_Generator_inst_2.count_dt\[0\]
+ _0580_ sky130_fd_sc_hd__a21oi_1
X_1066_ VPWR VGND VPWR VGND _0085_ _0445_ sky130_fd_sc_hd__inv_2
X_1135_ VGND VPWR _0517_ _0212_ _0208_ Signal_Generator_1_270phase_inst.count\[1\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_7_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ VGND VPWR VPWR VGND Signal_Generator_2_270phase_inst.count\[2\] _0396_ _0389_
+ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_9_Left_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 VGND VPWR Dead_Time_Generator_inst_1.dt\[4\] net30 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0704_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[0\] _0185_ Shift_Register_Inst.shift_state\[1\]
+ _0235_ _0183_ sky130_fd_sc_hd__or4b_1
X_0635_ VGND VPWR VPWR VGND _0187_ Dead_Time_Generator_inst_1.dt\[0\] _0186_ _0182_
+ sky130_fd_sc_hd__mux2_1
X_1118_ VPWR VGND VPWR VGND _0133_ _0442_ sky130_fd_sc_hd__inv_2
X_1049_ VPWR VGND VPWR VGND _0488_ net9 sky130_fd_sc_hd__inv_2
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Left_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0952_ VGND VPWR VPWR VGND _0419_ net6 Shift_Register_Inst.data_out\[13\] _0418_
+ sky130_fd_sc_hd__mux2_1
X_0883_ VGND VPWR _0370_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.count\[5\]
+ _0369_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_10_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1366_ Dead_Time_Generator_inst_3.count_dt\[3\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ net69 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1297_ VGND VPWR VPWR VGND clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0001_
+ _0080_ Signal_Generator_1_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1151_ VGND VPWR VGND VPWR Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0208_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0212_ _0533_ sky130_fd_sc_hd__mux4_1
X_1220_ VGND VPWR _0592_ net46 _0544_ _0591_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1082_ VPWR VGND VPWR VGND _0099_ _0498_ sky130_fd_sc_hd__inv_2
X_0866_ VPWR VGND Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] _0356_ Signal_Generator_2_90phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0935_ VPWR VGND Dead_Time_Generator_inst_1.clk _0407_ VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_0_23_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ VPWR VGND _0305_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
X_1349_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0046_
+ _0132_ Signal_Generator_2_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_0720_ VGND VPWR VGND VPWR _0244_ _0247_ _0246_ sky130_fd_sc_hd__or2b_1
X_0651_ VPWR VGND VGND VPWR Shift_Register_Inst.shift_state\[0\] _0196_ _0198_ sky130_fd_sc_hd__nor2_1
X_1134_ _0212_ Signal_Generator_1_90phase_inst.count\[1\] _0516_ _0208_ VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__and3b_1
X_1203_ VGND VPWR _0579_ _0577_ Dead_Time_Generator_inst_2.count_dt\[0\] _0578_ VPWR
+ VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Left_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1065_ VPWR VGND VPWR VGND _0084_ _0445_ sky130_fd_sc_hd__inv_2
X_0918_ VGND VPWR VPWR VGND Signal_Generator_2_270phase_inst.count\[2\] _0395_ _0392_
+ sky130_fd_sc_hd__xor2_1
X_0849_ VPWR VGND _0033_ _0327_ Signal_Generator_2_0phase_inst.direction Signal_Generator_2_0phase_inst.count\[4\]
+ _0343_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_38_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold6 net31 _0559_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0703_ VGND VPWR _0137_ _0234_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0634_ VPWR VGND VPWR VGND _0184_ _0185_ _0183_ _0186_ sky130_fd_sc_hd__or3_1
X_1117_ VPWR VGND VPWR VGND _0132_ _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1048_ VGND VPWR VGND VPWR Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[0\]
+ _0215_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[0\]
+ _0217_ _0487_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0882_ VGND VPWR _0369_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[3\]
+ _0368_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_27_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ VPWR VGND VPWR VGND _0418_ Dead_Time_Generator_inst_1.go sky130_fd_sc_hd__inv_2
XFILLER_0_10_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1365_ Dead_Time_Generator_inst_3.count_dt\[2\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0172_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1296_ VGND VPWR VPWR VGND clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0000_
+ _0079_ Signal_Generator_1_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1150_ VPWR VGND VGND VPWR _0532_ net41 _0409_ sky130_fd_sc_hd__or2_1
X_1081_ VPWR VGND VPWR VGND _0098_ _0498_ sky130_fd_sc_hd__inv_2
X_0865_ VPWR VGND VPWR VGND _0355_ _0346_ _0353_ _0051_ net71 sky130_fd_sc_hd__a22o_1
Xclkbuf_3_6__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR net27 clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
X_0934_ VGND VPWR VPWR VGND _0407_ Shift_Register_Inst.data_out\[14\] CLK_EXT CLK_PLL
+ sky130_fd_sc_hd__mux2_4
X_0796_ _0304_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0302_ _0303_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_1348_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0045_
+ _0131_ Signal_Generator_2_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1279_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0142_ _0063_ Shift_Register_Inst.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0650_ VPWR VGND VGND VPWR net79 _0197_ _0191_ _0153_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ VPWR VGND VPWR VGND _0083_ _0445_ sky130_fd_sc_hd__inv_2
X_1133_ _0208_ _0212_ _0515_ Signal_Generator_1_180phase_inst.count\[1\] VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__and3b_1
X_1202_ VGND VPWR VGND VPWR net30 _0578_ Dead_Time_Generator_inst_2.count_dt\[4\]
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0917_ VPWR VGND VPWR VGND _0394_ _0388_ _0393_ _0043_ Signal_Generator_2_270phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0779_ VGND VPWR VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0291_ _0284_
+ sky130_fd_sc_hd__xor2_1
X_0848_ _0343_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0323_ Signal_Generator_2_0phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xclkbuf_0_CLK_SR VGND VPWR VGND VPWR CLK_SR clknet_0_CLK_SR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold7 VGND VPWR net32 _0560_ VPWR VGND sky130_fd_sc_hd__buf_1
X_0633_ VPWR VGND VPWR VGND _0185_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ sky130_fd_sc_hd__or2_2
X_0702_ VGND VPWR VPWR VGND _0234_ Shift_Register_Inst.data_out\[15\] _0233_ net1
+ sky130_fd_sc_hd__mux2_1
X_1116_ VPWR VGND VPWR VGND _0131_ _0442_ sky130_fd_sc_hd__inv_2
X_1047_ VPWR VGND VGND VPWR net10 _0485_ _0486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0881_ VPWR VGND _0368_ Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[0\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_42_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ VGND VPWR net18 _0417_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1364_ Dead_Time_Generator_inst_3.count_dt\[1\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0171_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1295_ VPWR VGND VPWR VGND Signal_Generator_1_0phase_inst.direction _0078_ _0006_
+ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ VPWR VGND VPWR VGND _0097_ _0498_ sky130_fd_sc_hd__inv_2
X_0933_ VPWR VGND _0047_ _0390_ Signal_Generator_2_270phase_inst.direction Signal_Generator_2_270phase_inst.count\[4\]
+ _0406_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0864_ VPWR VGND VGND VPWR _0355_ _0349_ _0354_ sky130_fd_sc_hd__or2_1
X_0795_ VPWR VGND VPWR VGND _0303_ Signal_Generator_1_270phase_inst.direction sky130_fd_sc_hd__inv_2
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1347_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0044_
+ _0130_ Signal_Generator_2_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_1278_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0141_ _0062_ Shift_Register_Inst.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1201_ VPWR VGND VPWR VGND _0569_ net38 _0577_ _0574_ _0575_ _0576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1063_ VPWR VGND VPWR VGND _0082_ _0445_ sky130_fd_sc_hd__inv_2
X_1132_ VPWR VGND VPWR VGND _0512_ _0513_ _0510_ _0514_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0916_ VGND VPWR VGND VPWR _0391_ _0394_ _0393_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ VGND VPWR VPWR VGND Signal_Generator_1_180phase_inst.count\[2\] _0290_ _0287_
+ sky130_fd_sc_hd__xor2_1
X_0847_ VGND VPWR VPWR VGND _0032_ _0341_ _0340_ Signal_Generator_2_0phase_inst.direction
+ _0325_ _0342_ sky130_fd_sc_hd__a32o_1
Xhold8 net33 _0158_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0632_ VPWR VGND VGND VPWR _0184_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ sky130_fd_sc_hd__or2_1
X_0701_ VPWR VGND VGND VPWR _0233_ _0228_ _0191_ sky130_fd_sc_hd__or2_1
X_1115_ VPWR VGND VPWR VGND _0130_ _0442_ sky130_fd_sc_hd__inv_2
X_1046_ VGND VPWR VGND VPWR _0458_ _0481_ _0482_ _0483_ _0485_ _0484_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_45_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1029_ VGND VPWR VPWR VGND _0467_ _0465_ _0466_ _0468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_31_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ VGND VPWR VPWR VGND _0367_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0365_ _0366_ sky130_fd_sc_hd__o31a_2
XFILLER_0_12_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_42_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1363_ Dead_Time_Generator_inst_3.count_dt\[0\] clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
+ _0170_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1294_ Dead_Time_Generator_inst_4.go clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ _0157_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0932_ _0406_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0386_ Signal_Generator_2_270phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0863_ VGND VPWR VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0354_ _0347_
+ sky130_fd_sc_hd__xor2_1
X_0794_ VPWR VGND VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[0\]
+ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[3\]
+ _0302_ sky130_fd_sc_hd__or4_2
X_1346_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0043_
+ _0129_ Signal_Generator_2_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1277_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0140_ _0061_ Shift_Register_Inst.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1200_ _0576_ Dead_Time_Generator_inst_2.count_dt\[4\] net30 VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1062_ VPWR VGND VPWR VGND _0081_ _0445_ sky130_fd_sc_hd__inv_2
X_1131_ VPWR VGND VGND VPWR _0508_ _0509_ _0513_ sky130_fd_sc_hd__nor2_1
X_0915_ VPWR VGND VGND VPWR _0393_ _0392_ _0389_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0777_ VPWR VGND VPWR VGND _0289_ _0283_ _0288_ _0008_ net70 sky130_fd_sc_hd__a22o_1
X_0846_ VGND VPWR _0323_ _0342_ Signal_Generator_2_0phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0033_
+ _0112_ Signal_Generator_2_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_2
Xhold9 net34 Signal_Generator_1_90phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_29_Left_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0700_ VGND VPWR _0138_ _0232_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_0631_ VGND VPWR Shift_Register_Inst.shift_state\[4\] _0183_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_1114_ VPWR VGND VPWR VGND _0129_ _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1045_ VPWR VGND VPWR VGND _0217_ Signal_Generator_2_0phase_inst.count\[1\] _0215_
+ _0484_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0829_ VPWR VGND VPWR VGND _0028_ net54 sky130_fd_sc_hd__inv_2
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1028_ VPWR VGND _0467_ _0464_ net13 VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_26_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1293_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0156_ _0077_ Shift_Register_Inst.shift_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1362_ Dead_Time_Generator_inst_1.go clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
+ _0169_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0931_ VGND VPWR VPWR VGND _0046_ _0404_ _0403_ Signal_Generator_2_270phase_inst.direction
+ _0388_ _0405_ sky130_fd_sc_hd__a32o_1
X_0862_ VGND VPWR VPWR VGND Signal_Generator_2_90phase_inst.count\[2\] _0353_ _0350_
+ sky130_fd_sc_hd__xor2_1
X_0793_ VPWR VGND _0012_ _0285_ Signal_Generator_1_180phase_inst.direction Signal_Generator_1_180phase_inst.count\[4\]
+ _0301_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xrebuffer1 VPWR VGND VGND VPWR clknet_0_Dead_Time_Generator_inst_1.clk net26 sky130_fd_sc_hd__buf_8
X_1345_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0042_
+ _0128_ Signal_Generator_2_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1276_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0139_ _0060_ Shift_Register_Inst.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_1130_ VPWR VGND VPWR VGND _0507_ _0502_ _0501_ _0512_ sky130_fd_sc_hd__a21oi_1
X_1061_ VPWR VGND VPWR VGND _0080_ _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ VPWR VGND VGND VPWR Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ _0392_ sky130_fd_sc_hd__nor2_1
X_0845_ VPWR VGND VGND VPWR _0341_ Signal_Generator_2_0phase_inst.count\[4\] _0327_
+ sky130_fd_sc_hd__or2_1
X_0776_ VGND VPWR VGND VPWR _0286_ _0289_ _0288_ sky130_fd_sc_hd__or2b_1
X_1259_ VGND VPWR _0177_ _0621_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1328_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0032_
+ _0111_ Signal_Generator_2_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0630_ VPWR VGND _0182_ net1 VPWR VGND sky130_fd_sc_hd__buf_2
X_1044_ VGND VPWR _0483_ _0217_ _0215_ Signal_Generator_2_270phase_inst.count\[1\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_1113_ VPWR VGND VPWR VGND _0128_ _0442_ sky130_fd_sc_hd__inv_2
X_0759_ VPWR VGND VPWR VGND _0276_ _0262_ _0273_ _0024_ Signal_Generator_1_90phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_0828_ VPWR VGND VGND VPWR _0325_ _0328_ _0034_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Left_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ VPWR VGND _0466_ _0462_ net14 VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_Dead_Time_Generator_inst_1.clk VGND VPWR VGND VPWR net27 clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_14 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1361_ Dead_Time_Generator_inst_2.count_dt\[4\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ _0168_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1292_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0155_ _0076_ Shift_Register_Inst.shift_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0930_ VGND VPWR _0386_ _0405_ Signal_Generator_2_270phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_0861_ VPWR VGND VPWR VGND _0352_ _0346_ _0351_ _0050_ net71 sky130_fd_sc_hd__a22o_1
X_0792_ _0301_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0281_ Signal_Generator_1_180phase_inst.count\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xrebuffer2 VPWR VGND VPWR VGND net27 clknet_0_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1344_ VGND VPWR VPWR VGND clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0048_
+ _0127_ Signal_Generator_2_270phase_inst.direction sky130_fd_sc_hd__dfrtp_4
X_1275_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0138_ _0059_ Shift_Register_Inst.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1060_ VPWR VGND VPWR VGND _0079_ _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0913_ VPWR VGND VPWR VGND _0042_ net56 sky130_fd_sc_hd__inv_2
X_0775_ VPWR VGND VGND VPWR _0288_ _0287_ _0284_ sky130_fd_sc_hd__or2_1
X_0844_ VGND VPWR VPWR VGND Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0337_ _0340_ sky130_fd_sc_hd__or3b_1
X_1258_ VGND VPWR _0621_ _0594_ _0593_ _0620_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1327_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0031_
+ _0110_ Signal_Generator_2_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1189_ VPWR VGND VGND VPWR _0551_ _0563_ _0550_ _0568_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1112_ VPWR VGND VPWR VGND _0127_ _0442_ sky130_fd_sc_hd__inv_2
X_1043_ _0215_ _0217_ _0482_ Signal_Generator_2_180phase_inst.count\[1\] VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_43_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0827_ VGND VPWR _0328_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.count\[5\]
+ _0327_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0758_ VPWR VGND VPWR VGND _0275_ _0274_ _0265_ _0276_ sky130_fd_sc_hd__a21o_1
X_0689_ VGND VPWR VPWR VGND _0225_ Shift_Register_Inst.data_out\[11\] _0224_ net1
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1026_ VPWR VGND VGND VPWR net13 _0462_ net14 _0464_ _0465_ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ VGND VPWR VGND VPWR Dead_Time_Generator_inst_1.dt\[1\] _0448_ Dead_Time_Generator_inst_4.count_dt\[1\]
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1360_ Dead_Time_Generator_inst_2.count_dt\[3\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ _0167_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_1291_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0154_ _0075_ Shift_Register_Inst.shift_state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ VGND VPWR VGND VPWR _0349_ _0352_ _0351_ sky130_fd_sc_hd__or2b_1
X_0791_ VGND VPWR VPWR VGND _0011_ _0299_ _0298_ net74 _0283_ _0300_ sky130_fd_sc_hd__a32o_1
Xrebuffer3 VPWR VGND VPWR VGND net28 clknet_0_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dlygate4sd1_1
X_1343_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[5\] _0126_ _0040_
+ net29 sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1274_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0137_ _0058_ Shift_Register_Inst.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_0989_ VPWR VGND VPWR VGND _0062_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0912_ VPWR VGND VGND VPWR _0388_ _0391_ _0048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0774_ VPWR VGND VGND VPWR Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ _0287_ sky130_fd_sc_hd__nor2_1
X_0843_ VPWR VGND VPWR VGND _0339_ _0325_ _0336_ _0031_ Signal_Generator_2_0phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
X_1326_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0030_
+ _0109_ Signal_Generator_2_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_1188_ _0567_ Dead_Time_Generator_inst_1.count_dt\[1\] Dead_Time_Generator_inst_1.count_dt\[3\]
+ Dead_Time_Generator_inst_1.count_dt\[2\] net32 VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_1257_ VGND VPWR VPWR VGND Dead_Time_Generator_inst_4.count_dt\[1\] _0620_ _0616_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1111_ VPWR VGND VPWR VGND _0126_ _0442_ sky130_fd_sc_hd__inv_2
X_1042_ _0217_ Signal_Generator_2_90phase_inst.count\[1\] _0481_ _0215_ VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_9_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0757_ VPWR VGND _0275_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0688_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[2\] _0191_ _0188_ _0224_
+ sky130_fd_sc_hd__or3_1
X_0826_ VGND VPWR _0327_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ _0326_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1309_ VPWR VGND VPWR VGND Signal_Generator_1_180phase_inst.direction _0092_ _0013_
+ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1025_ VGND VPWR VGND VPWR _0457_ Signal_Generator_2_270phase_inst.count\[4\] _0458_
+ Signal_Generator_2_0phase_inst.count\[4\] _0464_ _0463_ sky130_fd_sc_hd__a221oi_2
X_0809_ VPWR VGND VPWR VGND _0313_ _0304_ _0311_ _0016_ Signal_Generator_1_270phase_inst.direction
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ VPWR VGND VPWR VGND _0447_ Dead_Time_Generator_inst_4.count_dt\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_37_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1290_ VGND VPWR VPWR VGND clknet_1_1__leaf_CLK_SR _0153_ _0074_ Shift_Register_Inst.shift_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_274 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer4 VPWR VGND VPWR VGND net29 clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
+ sky130_fd_sc_hd__dlygate4sd1_1
X_0790_ VGND VPWR _0281_ _0300_ Signal_Generator_1_180phase_inst.count\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_1342_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[4\] _0125_ _0039_
+ net29 sky130_fd_sc_hd__dfstp_2
X_1273_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0136_ _0057_ Shift_Register_Inst.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_0988_ VPWR VGND VPWR VGND _0061_ _0443_ sky130_fd_sc_hd__inv_2
X_0911_ VGND VPWR _0391_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.count\[5\]
+ _0390_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0842_ VPWR VGND VPWR VGND _0338_ _0337_ _0328_ _0339_ sky130_fd_sc_hd__a21o_1
X_0773_ VPWR VGND VPWR VGND _0007_ net57 sky130_fd_sc_hd__inv_2
X_1325_ VGND VPWR VPWR VGND clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0029_
+ _0108_ Signal_Generator_2_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1256_ VGND VPWR _0176_ _0619_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1187_ VPWR VGND VPWR VGND _0549_ _0545_ _0566_ _0160_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ VPWR VGND VPWR VGND _0125_ _0500_ sky130_fd_sc_hd__inv_2
X_1041_ VPWR VGND VPWR VGND _0476_ _0479_ _0478_ _0472_ _0480_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0825_ VPWR VGND _0326_ Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[0\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
X_0756_ VPWR VGND VPWR VGND _0274_ _0264_ sky130_fd_sc_hd__inv_2
X_0687_ VGND VPWR _0142_ _0223_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_1239_ VPWR VGND VGND VPWR Dead_Time_Generator_inst_3.count_dt\[1\] _0608_ _0605_
+ sky130_fd_sc_hd__nand2_1
X_1308_ VGND VPWR VPWR VGND clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0026_
+ _0091_ Signal_Generator_1_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Left_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1024_ VPWR VGND VPWR VGND _0460_ Signal_Generator_2_180phase_inst.count\[4\] _0459_
+ _0463_ Signal_Generator_2_90phase_inst.count\[4\] sky130_fd_sc_hd__a22o_1
X_0808_ VPWR VGND VGND VPWR _0313_ _0307_ _0312_ sky130_fd_sc_hd__or2_1
X_0739_ VPWR VGND VPWR VGND _0261_ Signal_Generator_1_90phase_inst.direction sky130_fd_sc_hd__inv_2
XFILLER_0_22_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ VPWR VGND VPWR VGND _0446_ Dead_Time_Generator_inst_4.count_dt\[3\] sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_CLK_SR VGND VPWR VGND VPWR clknet_0_CLK_SR clknet_1_0__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Left_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1341_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[3\] _0124_ _0038_
+ net29 sky130_fd_sc_hd__dfstp_1
X_1272_ VGND VPWR VPWR VGND clknet_1_0__leaf_CLK_SR _0135_ _0056_ Shift_Register_Inst.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_0987_ VPWR VGND VPWR VGND _0060_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0910_ VGND VPWR _0390_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ _0389_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0772_ VPWR VGND VGND VPWR _0283_ _0286_ _0013_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0841_ VPWR VGND _0338_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1186_ VGND VPWR _0563_ _0566_ _0551_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_1255_ VGND VPWR _0619_ _0594_ _0593_ _0618_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1324_ VGND VPWR VPWR VGND clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0028_
+ _0107_ Signal_Generator_2_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1040_ VGND VPWR _0479_ _0474_ net11 _0475_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0824_ VGND VPWR VPWR VGND _0325_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0323_ _0324_ sky130_fd_sc_hd__o31a_2
X_0755_ VPWR VGND VGND VPWR _0260_ _0273_ _0272_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Left_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0686_ VGND VPWR VPWR VGND _0223_ Shift_Register_Inst.data_out\[10\] _0222_ net1
+ sky130_fd_sc_hd__mux2_1
X_1307_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[4\] _0090_ _0025_
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1169_ VPWR VGND VPWR VGND _0551_ net52 sky130_fd_sc_hd__inv_2
X_1238_ VPWR VGND VPWR VGND _0170_ _0607_ _0605_ _0593_ _0594_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_42_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1023_ VGND VPWR VGND VPWR _0457_ Signal_Generator_2_270phase_inst.count\[5\] _0458_
+ Signal_Generator_2_0phase_inst.count\[5\] _0462_ _0461_ sky130_fd_sc_hd__a221oi_2
X_0738_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[0\]
+ Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[3\]
+ _0260_ sky130_fd_sc_hd__or4_2
X_0807_ VGND VPWR VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] _0312_ _0305_
+ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0669_ VGND VPWR VPWR VGND _0211_ _0208_ _0210_ _0182_ sky130_fd_sc_hd__mux2_1
Xhold50 net75 Dead_Time_Generator_inst_3.count_dt\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ VPWR VGND VPWR VGND _0077_ _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_243 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1340_ VPWR VGND VPWR VGND Signal_Generator_2_180phase_inst.count\[2\] _0123_ _0037_
+ net29 sky130_fd_sc_hd__dfstp_2
XFILLER_0_23_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1271_ VPWR VGND VPWR VGND _0594_ _0593_ _0606_ _0181_ sky130_fd_sc_hd__a21oi_1
X_0986_ VPWR VGND VPWR VGND _0059_ _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0840_ VPWR VGND VPWR VGND _0337_ _0327_ sky130_fd_sc_hd__inv_2
X_0771_ VGND VPWR _0286_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.count\[5\]
+ _0285_ VPWR VGND sky130_fd_sc_hd__and3_1
X_1323_ VPWR VGND VPWR VGND Signal_Generator_2_0phase_inst.direction _0106_ _0034_
+ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_2
X_1254_ VPWR VGND VGND VPWR _0616_ _0617_ _0618_ sky130_fd_sc_hd__nor2_1
X_1185_ VPWR VGND VPWR VGND _0549_ _0545_ _0565_ _0159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ VPWR VGND _0431_ Shift_Register_Inst.data_out\[10\] Shift_Register_Inst.data_out\[9\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0754_ VPWR VGND Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] _0272_ Signal_Generator_1_90phase_inst.count\[3\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0685_ VPWR VGND VPWR VGND Shift_Register_Inst.shift_state\[2\] _0201_ _0188_ _0222_
+ sky130_fd_sc_hd__or3_1
X_0823_ VPWR VGND VPWR VGND _0324_ Signal_Generator_2_0phase_inst.direction sky130_fd_sc_hd__inv_2
X_1306_ VPWR VGND VPWR VGND Signal_Generator_1_90phase_inst.count\[3\] _0089_ _0024_
+ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__dfstp_1
XFILLER_0_19_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ VPWR VGND VPWR VGND _0115_ _0499_ sky130_fd_sc_hd__inv_2
X_1168_ VPWR VGND VPWR VGND _0550_ net50 sky130_fd_sc_hd__inv_2
X_1237_ VPWR VGND VGND VPWR net62 _0606_ _0607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ VPWR VGND VPWR VGND _0460_ Signal_Generator_2_180phase_inst.count\[5\] _0459_
+ _0461_ Signal_Generator_2_90phase_inst.count\[5\] sky130_fd_sc_hd__a22o_1
X_0737_ VPWR VGND _0005_ _0243_ Signal_Generator_1_0phase_inst.direction Signal_Generator_1_0phase_inst.count\[4\]
+ _0259_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0668_ VPWR VGND VGND VPWR _0210_ _0193_ _0209_ sky130_fd_sc_hd__or2_1
X_0806_ VGND VPWR VPWR VGND Signal_Generator_1_270phase_inst.count\[2\] _0311_ _0308_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold40 VGND VPWR Signal_Generator_2_180phase_inst.count\[0\] net65 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold51 net76 Shift_Register_Inst.shift_state\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1005_ VPWR VGND VPWR VGND _0076_ _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
.ends

