magic
tech sky130A
timestamp 1698344643
<< checkpaint >>
rect -630 56970 37830 133430
rect -630 -630 29030 56970
<< metal2 >>
rect 3000 127060 5200 127600
rect 3000 126870 4960 127060
rect 3000 126000 5200 126870
rect 3000 62560 5740 62800
rect 5930 62560 6800 62800
rect 3000 61200 6800 62560
rect 3000 52240 6800 53600
rect 3000 52000 5740 52240
rect 5930 52000 6800 52240
rect 3000 5749 4962 6000
rect 3000 5200 5300 5749
<< metal3 >>
rect 6000 128600 36000 131600
rect 1000 99600 4000 125600
rect 33000 101600 36000 128600
rect 1000 90600 31000 99600
rect 1000 63600 4000 90600
rect 33000 61600 36000 88600
rect 6000 58600 36000 61600
rect 6000 53600 27800 58600
rect 1000 32800 4000 51600
rect 24800 34800 27800 53600
rect 1000 24800 22800 32800
rect 1000 7000 4000 24800
rect 24800 4000 27800 22800
rect 6000 1000 27800 4000
<< metal4 >>
rect 6000 128600 36000 131600
rect 1000 99600 4000 125600
rect 33000 101600 36000 128600
rect 1000 90600 31000 99600
rect 1000 63600 4000 90600
rect 33000 61600 36000 88600
rect 6000 58600 36000 61600
rect 6000 53600 27800 58600
rect 1000 32800 4000 51600
rect 24800 34800 27800 53600
rect 1000 24800 22800 32800
rect 1000 7000 4000 24800
rect 24800 4000 27800 22800
rect 6000 1000 27800 4000
<< metal5 >>
rect 6000 128600 36000 131600
rect 1000 99600 4000 125600
rect 33000 101600 36000 128600
rect 1000 90600 31000 99600
rect 1000 63600 4000 90600
rect 33000 61600 36000 88600
rect 6000 58600 36000 61600
rect 6000 53600 27800 58600
rect 1000 32800 4000 51600
rect 24800 34800 27800 53600
rect 1000 24800 22800 32800
rect 1000 7000 4000 24800
rect 24800 4000 27800 22800
rect 6000 1000 27800 4000
use nmos_waffle_32x32  nmos_waffle_32x32_0
timestamp 1698344533
transform 1 0 5925 0 1 5975
box -5925 -5975 22475 22425
use nmos_waffle_32x32  nmos_waffle_32x32_1
timestamp 1698344533
transform 0 1 5975 -1 0 51275
box -5925 -5975 22475 22425
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1684343764
transform 0 1 5975 1 0 63525
box -5925 -5975 31275 31225
use pmos_waffle_48x48  pmos_waffle_48x48_1
timestamp 1684343764
transform 1 0 5925 0 -1 126825
box -5925 -5975 31275 31225
<< labels >>
rlabel metal5 6000 129600 7000 130600 7 VP
rlabel metal2 3000 126600 4000 127600 7 s1
rlabel metal5 1000 94600 2000 95600 7 fc1
rlabel metal2 3000 61600 4000 62600 7 s2
rlabel metal5 6000 56600 22400 57600 7 out
rlabel metal2 3000 52600 4000 53600 7 s3
rlabel metal5 1000 28300 2000 29300 7 fc2
rlabel metal2 3000 5500 4000 6000 7 s4
rlabel metal5 6000 2000 7000 3000 7 VN
<< end >>
