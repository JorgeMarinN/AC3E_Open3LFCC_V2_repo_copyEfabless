magic
tech sky130A
timestamp 1698343393
<< checkpaint >>
rect -6555 -6605 28605 28555
<< nwell >>
rect -1125 22000 0 23125
rect 22000 22000 23175 23125
rect -1125 -1175 0 0
rect 22000 -1175 23175 0
<< pwell >>
rect -5925 23125 27975 27925
rect -5925 -1175 -1125 23125
rect 23175 -1175 27975 23125
rect -5925 -5975 27975 -1175
<< mvpmos >>
rect 22000 22031 22050 22469
rect -469 -50 -31 0
rect 22081 -50 22519 0
rect 22000 -519 22050 -81
<< mvpdiff >>
rect 22079 22469 22521 22471
rect -29 22463 0 22469
rect -29 22064 -23 22463
rect -64 22037 -23 22064
rect -6 22037 0 22463
rect -64 22031 0 22037
rect 21997 22031 22000 22469
rect 22050 22463 22521 22469
rect 22050 22037 22056 22463
rect 22073 22415 22521 22463
rect 22073 22085 22135 22415
rect 22465 22085 22521 22415
rect 22073 22037 22521 22085
rect 22050 22031 22521 22037
rect -64 22029 -31 22031
rect -469 22023 -31 22029
rect -469 22006 -463 22023
rect -37 22006 -31 22023
rect -469 22000 -31 22006
rect 22079 22029 22521 22031
rect 22081 22023 22519 22029
rect 22081 22006 22087 22023
rect 22513 22006 22519 22023
rect 22081 22000 22519 22006
rect -469 0 -31 3
rect 22081 0 22519 3
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 22081 -56 22519 -50
rect 22081 -73 22087 -56
rect 22513 -73 22519 -56
rect 22081 -79 22519 -73
rect 22081 -81 22114 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 21997 -519 22000 -81
rect 22050 -87 22114 -81
rect 22050 -513 22056 -87
rect 22073 -114 22114 -87
rect 22073 -513 22079 -114
rect 22050 -519 22079 -513
rect -471 -521 -29 -519
<< mvpdiffc >>
rect -23 22037 -6 22463
rect 22056 22037 22073 22463
rect -463 22006 -37 22023
rect 22087 22006 22513 22023
rect -463 -73 -37 -56
rect 22087 -73 22513 -56
rect -23 -513 -6 -87
rect 22056 -513 22073 -87
<< mvpsubdiff >>
rect -5525 27513 27575 27525
rect -5525 -5563 -5513 27513
rect -1537 23525 23587 23537
rect -1537 -1575 -1525 23525
rect 23575 -1575 23587 23525
rect -1537 -1587 23587 -1575
rect 27563 -5563 27575 27513
rect -5525 -5575 27575 -5563
<< mvnsubdiff >>
rect -1025 23013 0 23025
rect -1025 22017 -1013 23013
rect -17 22737 0 23013
rect -737 22725 0 22737
rect 22000 23013 23075 23025
rect 22000 22725 22787 22737
rect -737 22017 -725 22725
rect -1025 22000 -725 22017
rect 22135 22403 22465 22415
rect 22135 22097 22147 22403
rect 22453 22097 22465 22403
rect 22135 22085 22465 22097
rect 22775 22017 22787 22725
rect 23063 22017 23075 23013
rect 22775 22000 23075 22017
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 22775 -775 22787 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 22000 -787 22787 -775
rect 23063 -1063 23075 0
rect 22000 -1075 23075 -1063
<< mvpsubdiffcont >>
rect -5513 23537 27563 27513
rect -5513 -1587 -1537 23537
rect 23587 -1587 27563 23537
rect -5513 -5563 27563 -1587
<< mvnsubdiffcont >>
rect -1013 22737 -17 23013
rect -1013 22017 -737 22737
rect 22000 22737 23063 23013
rect 22147 22097 22453 22403
rect 22787 22017 23063 22737
rect -1013 -787 -737 0
rect -403 -453 -97 -147
rect -1013 -1063 -17 -787
rect 22787 -787 23063 0
rect 22000 -1063 23063 -787
<< poly >>
rect -550 22542 0 22550
rect -550 22508 -542 22542
rect -508 22508 0 22542
rect -550 22500 0 22508
rect 22000 22542 22600 22550
rect 22000 22508 22008 22542
rect 22042 22508 22558 22542
rect 22592 22508 22600 22542
rect 22000 22500 22600 22508
rect -550 22000 -500 22500
rect 22000 22469 22050 22500
rect 22000 22000 22050 22031
rect 22550 22000 22600 22500
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -50 0 0
rect 22000 -8 22081 0
rect 22000 -42 22008 -8
rect 22042 -42 22081 -8
rect 22000 -50 22081 -42
rect 22519 -8 22600 0
rect 22519 -42 22558 -8
rect 22592 -42 22600 -8
rect 22519 -50 22600 -42
rect -550 -550 -500 -50
rect 22000 -81 22050 -50
rect 22000 -550 22050 -519
rect 22550 -550 22600 -50
rect -550 -558 0 -550
rect -550 -592 -542 -558
rect -508 -592 0 -558
rect -550 -600 0 -592
rect 22000 -558 22600 -550
rect 22000 -592 22008 -558
rect 22042 -592 22558 -558
rect 22592 -592 22600 -558
rect 22000 -600 22600 -592
<< polycont >>
rect -542 22508 -508 22542
rect 22008 22508 22042 22542
rect 22558 22508 22592 22542
rect -542 -42 -508 -8
rect 22008 -42 22042 -8
rect 22558 -42 22592 -8
rect -542 -592 -508 -558
rect 22008 -592 22042 -558
rect 22558 -592 22592 -558
<< locali >>
rect -5525 27513 27575 27525
rect -5525 -5563 -5513 27513
rect -1537 23525 23587 23537
rect -1537 -1575 -1525 23525
rect -1025 23013 0 23025
rect -1025 22017 -1013 23013
rect -17 22737 0 23013
rect -737 22725 0 22737
rect 22000 23013 23075 23025
rect 22000 22725 22787 22737
rect -737 22017 -725 22725
rect -550 22542 -500 22550
rect -550 22508 -542 22542
rect -508 22508 -500 22542
rect -550 22500 -500 22508
rect 22000 22542 22050 22550
rect 22000 22508 22008 22542
rect 22042 22508 22050 22542
rect 22000 22500 22050 22508
rect 22550 22542 22600 22550
rect 22550 22508 22558 22542
rect 22592 22508 22600 22542
rect 22550 22500 22600 22508
rect 22073 22471 22527 22477
rect -23 22463 -6 22471
rect -64 22037 -23 22064
rect -64 22029 -6 22037
rect 22056 22463 22527 22471
rect 22073 22415 22527 22463
rect 22073 22085 22135 22415
rect 22465 22085 22527 22415
rect 22073 22037 22527 22085
rect 22056 22029 22527 22037
rect -64 22023 -29 22029
rect 22073 22023 22527 22029
rect -1025 22000 -725 22017
rect -471 22006 -463 22023
rect -37 22006 -29 22023
rect 22079 22006 22087 22023
rect 22513 22006 22521 22023
rect 22775 22017 22787 22725
rect 23063 22017 23075 23013
rect 22775 22000 23075 22017
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 22000 -8 22050 0
rect 22000 -42 22008 -8
rect 22042 -42 22050 -8
rect 22000 -50 22050 -42
rect 22550 -8 22600 0
rect 22550 -42 22558 -8
rect 22592 -42 22600 -8
rect 22550 -50 22600 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 22079 -73 22087 -56
rect 22513 -73 22521 -56
rect -477 -79 -23 -73
rect 22079 -79 22114 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 22056 -87 22114 -79
rect 22073 -114 22114 -87
rect 22056 -521 22073 -513
rect -477 -527 -23 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 22000 -558 22050 -550
rect 22000 -592 22008 -558
rect 22042 -592 22050 -558
rect 22000 -600 22050 -592
rect 22550 -558 22600 -550
rect 22550 -592 22558 -558
rect 22592 -592 22600 -558
rect 22550 -600 22600 -592
rect 22775 -775 22787 0
rect -737 -787 0 -775
rect -17 -1063 0 -787
rect -1025 -1075 0 -1063
rect 22000 -787 22787 -775
rect 23063 -1063 23075 0
rect 22000 -1075 23075 -1063
rect 23575 -1575 23587 23525
rect -1537 -1587 23587 -1575
rect 27563 -5563 27575 27513
rect -5525 -5575 27575 -5563
<< viali >>
rect -5513 23537 27563 27513
rect -5513 -1587 -1537 23537
rect -1013 22737 -19 23013
rect -1013 22019 -737 22737
rect 22000 22737 23063 23013
rect -542 22508 -508 22542
rect 22008 22508 22042 22542
rect 22558 22508 22592 22542
rect -23 22037 -6 22463
rect 22056 22037 22073 22463
rect 22135 22403 22465 22415
rect 22135 22097 22147 22403
rect 22147 22097 22453 22403
rect 22453 22097 22465 22403
rect 22135 22085 22465 22097
rect -463 22006 -37 22023
rect 22087 22006 22513 22023
rect 22787 22019 23063 22737
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 22008 -42 22042 -8
rect 22558 -42 22592 -8
rect -463 -73 -37 -56
rect 22087 -73 22513 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 22056 -513 22073 -87
rect -542 -592 -508 -558
rect 22008 -592 22042 -558
rect 22558 -592 22592 -558
rect -1013 -1063 -19 -787
rect 22787 -787 23063 0
rect 22000 -1063 23063 -787
rect 23587 -1587 27563 23537
rect -5513 -5563 27563 -1587
<< metal1 >>
rect -5525 27513 27575 27525
rect -5525 -5563 -5513 27513
rect -1537 23525 23587 23537
rect -1537 -1575 -1525 23525
rect -1025 23013 0 23025
rect -1025 22019 -1013 23013
rect -19 22737 0 23013
rect -737 22725 0 22737
rect 22000 23013 23075 23025
rect 22000 22725 22787 22737
rect -737 22019 -725 22725
rect -550 22542 -500 22550
rect -550 22508 -542 22542
rect -508 22508 -500 22542
rect -550 22500 -500 22508
rect 22000 22542 22050 22550
rect 22000 22508 22008 22542
rect 22042 22508 22050 22542
rect 22000 22500 22050 22508
rect 22550 22542 22600 22550
rect 22550 22508 22558 22542
rect 22592 22508 22600 22542
rect 22550 22500 22600 22508
rect -474 22469 -26 22474
rect 22076 22469 22524 22474
rect -474 22463 -3 22469
rect -474 22415 -23 22463
rect -474 22085 -415 22415
rect -85 22085 -23 22415
rect -474 22037 -23 22085
rect -6 22037 -3 22463
rect -474 22031 -3 22037
rect 22053 22463 22524 22469
rect 22053 22037 22056 22463
rect 22073 22415 22524 22463
rect 22073 22085 22135 22415
rect 22465 22085 22524 22415
rect 22073 22037 22524 22085
rect 22053 22031 22524 22037
rect -474 22026 -26 22031
rect 22076 22026 22524 22031
rect -1025 22000 -725 22019
rect -469 22023 -31 22026
rect -469 22006 -463 22023
rect -37 22006 -31 22023
rect -469 22003 -31 22006
rect 22081 22023 22519 22026
rect 22081 22006 22087 22023
rect 22513 22006 22519 22023
rect 22081 22003 22519 22006
rect 22775 22019 22787 22725
rect 23063 22019 23075 23013
rect 22775 22000 23075 22019
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 22000 -8 22050 0
rect 22000 -42 22008 -8
rect 22042 -42 22050 -8
rect 22000 -50 22050 -42
rect 22550 -8 22600 0
rect 22550 -42 22558 -8
rect 22592 -42 22600 -8
rect 22550 -50 22600 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 22081 -56 22519 -53
rect 22081 -73 22087 -56
rect 22513 -73 22519 -56
rect 22081 -76 22519 -73
rect -474 -81 -26 -76
rect 22076 -81 22524 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 22053 -87 22524 -81
rect 22053 -513 22056 -87
rect 22073 -135 22524 -87
rect 22073 -465 22135 -135
rect 22465 -465 22524 -135
rect 22073 -513 22524 -465
rect 22053 -519 22524 -513
rect -474 -524 -26 -519
rect 22076 -524 22524 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 22000 -558 22050 -550
rect 22000 -592 22008 -558
rect 22042 -592 22050 -558
rect 22000 -600 22050 -592
rect 22550 -558 22600 -550
rect 22550 -592 22558 -558
rect 22592 -592 22600 -558
rect 22550 -600 22600 -592
rect 22775 -775 22787 0
rect -737 -787 0 -775
rect -19 -1063 0 -787
rect -1025 -1075 0 -1063
rect 22000 -787 22787 -775
rect 23063 -1063 23075 0
rect 22000 -1075 23075 -1063
rect 23575 -1575 23587 23525
rect -1537 -1587 23587 -1575
rect 27563 -5563 27575 27513
rect -5525 -5575 27575 -5563
<< via1 >>
rect -5513 23537 27563 27513
rect -5513 1117 -1537 23525
rect 22088 22825 22188 22925
rect -542 22508 -508 22542
rect 22008 22508 22042 22542
rect 22558 22508 22592 22542
rect -415 22085 -85 22415
rect 22135 22085 22465 22415
rect 22875 22038 22975 22138
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 22008 -42 22042 -8
rect 22558 -42 22592 -8
rect -415 -465 -85 -135
rect 22135 -465 22465 -135
rect -542 -592 -508 -558
rect 22008 -592 22042 -558
rect 22558 -592 22592 -558
rect -138 -975 -38 -875
rect 23587 -1587 27563 23537
rect -495 -5563 27563 -1587
<< metal2 >>
rect -5525 27513 27575 27525
rect -5525 23537 -5513 27513
rect -5525 23525 23587 23537
rect -5525 1117 -5513 23525
rect -1537 1117 -1525 23525
rect 22078 22925 22198 22935
rect 22078 22825 22088 22925
rect 22188 22825 22198 22925
rect 22078 22815 22198 22825
rect -725 22542 0 22725
rect -725 22508 -542 22542
rect -508 22508 0 22542
rect -725 22500 0 22508
rect 22000 22542 22775 22725
rect 22000 22508 22008 22542
rect 22042 22508 22558 22542
rect 22592 22508 22775 22542
rect 22000 22500 22775 22508
rect -725 22000 -500 22500
rect -425 22415 -75 22425
rect -425 22085 -415 22415
rect -85 22085 -75 22415
rect -425 22075 -75 22085
rect 22000 22000 22050 22500
rect 22125 22415 22475 22425
rect 22125 22085 22135 22415
rect 22465 22085 22475 22415
rect 22125 22075 22475 22085
rect 22550 22000 22775 22500
rect 22865 22138 22985 22148
rect 22865 22038 22875 22138
rect 22975 22038 22985 22138
rect 22865 22028 22985 22038
rect -725 -8 0 0
rect -725 -42 -542 -8
rect -508 -42 0 -8
rect -725 -50 0 -42
rect 22000 -8 22775 0
rect 22000 -42 22008 -8
rect 22042 -42 22558 -8
rect 22592 -42 22775 -8
rect 22000 -50 22775 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 22000 -550 22050 -50
rect 22125 -135 22475 -125
rect 22125 -465 22135 -135
rect 22465 -465 22475 -135
rect 22125 -475 22475 -465
rect 22550 -550 22775 -50
rect -725 -558 0 -550
rect -725 -592 -542 -558
rect -508 -592 0 -558
rect -725 -775 0 -592
rect 22000 -558 22775 -550
rect 22000 -592 22008 -558
rect 22042 -592 22558 -558
rect 22592 -592 22775 -558
rect 22000 -775 22775 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 23575 -1575 23587 23525
rect -507 -1587 23587 -1575
rect -507 -5563 -495 -1587
rect 27563 -5563 27575 27513
rect -507 -5575 27575 -5563
<< via2 >>
rect 22088 22825 22188 22925
rect -310 22190 -190 22310
rect 22240 22190 22360 22310
rect 22875 22038 22975 22138
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 22240 -360 22360 -240
rect -138 -975 -38 -875
<< metal3 >>
rect -2525 23525 22575 24525
rect -2525 22638 -1525 23525
rect -638 22638 -186 23525
rect -2525 22314 -186 22638
rect -88 22412 0 23025
tri -186 22314 -88 22412 sw
tri -88 22324 0 22412 ne
rect 22000 22925 22364 23025
rect 22000 22825 22088 22925
rect 22188 22825 22364 22925
rect 22000 22324 22364 22825
rect -2525 22310 -88 22314
rect -2525 22190 -310 22310
rect -190 22226 -88 22310
tri -88 22226 0 22314 sw
rect -190 22190 0 22226
rect -2525 22186 0 22190
rect -2525 -575 -1525 22186
tri -412 22088 -314 22186 ne
rect -314 22088 0 22186
rect -1025 22000 -412 22088
tri -412 22000 -324 22088 sw
tri -314 22000 -226 22088 ne
rect -226 22000 0 22088
tri 22000 22226 22098 22324 ne
rect 22098 22314 22364 22324
tri 22364 22314 22462 22412 sw
rect 23575 22314 24575 22525
rect 22098 22310 24575 22314
rect 22098 22226 22240 22310
tri 22000 22138 22088 22226 sw
tri 22098 22138 22186 22226 ne
rect 22186 22190 22240 22226
rect 22360 22190 24575 22310
rect 22186 22138 24575 22190
rect 22000 22058 22088 22138
tri 22088 22058 22168 22138 sw
tri 22186 22058 22266 22138 ne
rect 22266 22058 22875 22138
rect 22000 22000 22168 22058
tri 22168 22000 22226 22058 sw
tri 22266 22000 22324 22058 ne
rect 22324 22038 22875 22058
rect 22975 22038 24575 22138
rect 22324 22000 24575 22038
rect 23575 0 24575 22000
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 22000 -40 22226 0
tri 22226 -40 22266 0 sw
tri 22324 -40 22364 0 ne
rect 22364 -40 24575 0
rect 22000 -138 22266 -40
tri 22266 -138 22364 -40 sw
tri 22364 -138 22462 -40 ne
rect 22462 -138 24575 -40
rect 22000 -226 22364 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 22000 -324 22098 -226 ne
rect 22098 -236 22364 -226
tri 22364 -236 22462 -138 sw
rect 22098 -240 23075 -236
rect 22098 -324 22240 -240
tri 22000 -364 22040 -324 sw
tri 22098 -364 22138 -324 ne
rect 22138 -360 22240 -324
rect 22360 -360 23075 -240
rect 22138 -364 23075 -360
rect 22000 -462 22040 -364
tri 22040 -462 22138 -364 sw
tri 22138 -462 22236 -364 ne
rect 22000 -1575 22138 -462
rect 22236 -688 23075 -364
rect 22236 -1075 22688 -688
rect 23575 -1575 24575 -138
rect -525 -2575 24575 -1575
<< via3 >>
rect 22088 22825 22188 22925
rect -310 22190 -190 22310
rect 22240 22190 22360 22310
rect 22875 22038 22975 22138
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect -138 -975 -38 -875
rect 22240 -360 22360 -240
<< metal4 >>
rect -2525 23525 22575 24525
rect -2525 22638 -1525 23525
rect -638 22638 -186 23525
rect -2525 22314 -186 22638
rect -88 22412 0 23025
tri -186 22314 -88 22412 sw
tri -88 22324 0 22412 ne
rect 22000 22925 22364 23025
rect 22000 22825 22088 22925
rect 22188 22825 22364 22925
rect 22000 22324 22364 22825
rect -2525 22310 -88 22314
rect -2525 22190 -310 22310
rect -190 22226 -88 22310
tri -88 22226 0 22314 sw
rect -190 22190 0 22226
rect -2525 22186 0 22190
rect -2525 -575 -1525 22186
tri -412 22088 -314 22186 ne
rect -314 22088 0 22186
rect -1025 22000 -412 22088
tri -412 22000 -324 22088 sw
tri -314 22000 -226 22088 ne
rect -226 22000 0 22088
tri 22000 22226 22098 22324 ne
rect 22098 22314 22364 22324
tri 22364 22314 22462 22412 sw
rect 23575 22314 24575 22525
rect 22098 22310 24575 22314
rect 22098 22226 22240 22310
tri 22000 22138 22088 22226 sw
tri 22098 22138 22186 22226 ne
rect 22186 22190 22240 22226
rect 22360 22190 24575 22310
rect 22186 22138 24575 22190
rect 22000 22058 22088 22138
tri 22088 22058 22168 22138 sw
tri 22186 22058 22266 22138 ne
rect 22266 22058 22875 22138
rect 22000 22000 22168 22058
tri 22168 22000 22226 22058 sw
tri 22266 22000 22324 22058 ne
rect 22324 22038 22875 22058
rect 22975 22038 24575 22138
rect 22324 22000 24575 22038
rect 23575 0 24575 22000
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 0 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -138 0 -40
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -226 0 -138 ne
rect 22000 -40 22226 0
tri 22226 -40 22266 0 sw
tri 22324 -40 22364 0 ne
rect 22364 -40 24575 0
rect 22000 -138 22266 -40
tri 22266 -138 22364 -40 sw
tri 22364 -138 22462 -40 ne
rect 22462 -138 24575 -40
rect 22000 -226 22364 -138
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri -412 -462 -314 -364 ne
rect -314 -875 0 -364
rect -314 -975 -138 -875
rect -38 -975 0 -875
rect -314 -1575 0 -975
tri 22000 -324 22098 -226 ne
rect 22098 -236 22364 -226
tri 22364 -236 22462 -138 sw
rect 22098 -240 23075 -236
rect 22098 -324 22240 -240
tri 22000 -364 22040 -324 sw
tri 22098 -364 22138 -324 ne
rect 22138 -360 22240 -324
rect 22360 -360 23075 -240
rect 22138 -364 23075 -360
rect 22000 -462 22040 -364
tri 22040 -462 22138 -364 sw
tri 22138 -462 22236 -364 ne
rect 22000 -1575 22138 -462
rect 22236 -688 23075 -364
rect 22236 -1075 22688 -688
rect 23575 -1575 24575 -138
rect -525 -2575 24575 -1575
<< via4 >>
rect -310 22190 -190 22310
rect 22240 22190 22360 22310
rect -310 -360 -190 -240
rect 22240 -360 22360 -240
<< metal5 >>
rect -2525 23525 22575 24525
rect -2525 22603 -1525 23525
rect -603 22603 -292 23525
rect -2525 22310 -292 22603
tri -292 22310 -154 22448 sw
rect -53 22447 0 23025
tri -53 22394 0 22447 ne
rect 22000 22394 22258 23025
rect -2525 22292 -310 22310
rect -2525 -575 -1525 22292
tri -448 22156 -312 22292 ne
rect -312 22190 -310 22292
rect -190 22190 -154 22310
rect -312 22156 -154 22190
tri -154 22156 0 22310 sw
rect -1025 22000 -447 22053
tri -447 22000 -394 22053 sw
tri -312 22000 -156 22156 ne
rect -156 22000 0 22156
tri 22000 22156 22238 22394 ne
rect 22238 22310 22258 22394
tri 22258 22310 22396 22448 sw
rect 22238 22190 22240 22310
rect 22360 22208 22396 22310
tri 22396 22208 22498 22310 sw
rect 23575 22208 24575 22525
rect 22360 22190 24575 22208
rect 22238 22156 24575 22190
tri 22000 22000 22156 22156 sw
tri 22238 22000 22394 22156 ne
rect 22394 22000 24575 22156
rect 23575 0 24575 22000
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 0 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -156 0 -103 ne
rect 22000 -103 22156 0
tri 22156 -103 22259 0 sw
tri 22394 -103 22497 0 ne
rect 22497 -103 24575 0
rect 22000 -156 22259 -103
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
rect -208 -1575 0 -394
tri 22000 -394 22238 -156 ne
rect 22238 -240 22259 -156
tri 22259 -240 22396 -103 sw
rect 22238 -360 22240 -240
rect 22360 -342 22396 -240
tri 22396 -342 22498 -240 sw
rect 22360 -360 23075 -342
rect 22238 -394 23075 -360
tri 22000 -497 22103 -394 sw
rect 22000 -1575 22103 -497
tri 22238 -498 22342 -394 ne
rect 22342 -653 23075 -394
rect 22342 -1075 22653 -653
rect 23575 -1575 24575 -103
rect -525 -2575 24575 -1575
use pmos_drain_frame_lt  pmos_drain_frame_lt_0 waffle_cells
timestamp 1675433017
transform 1 0 -550 0 1 0
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_1
timestamp 1675433017
transform 0 -1 1100 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_2
timestamp 1675433017
transform 1 0 -550 0 1 1100
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_3
timestamp 1675433017
transform 0 -1 2200 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_4
timestamp 1675433017
transform 1 0 -550 0 1 2200
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_5
timestamp 1675433017
transform 0 -1 3300 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_6
timestamp 1675433017
transform 1 0 -550 0 1 3300
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_7
timestamp 1675433017
transform 0 -1 4400 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_8
timestamp 1675433017
transform 1 0 -550 0 1 4400
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_9
timestamp 1675433017
transform 0 -1 5500 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_10
timestamp 1675433017
transform 1 0 -550 0 1 5500
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_11
timestamp 1675433017
transform 0 -1 6600 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_12
timestamp 1675433017
transform 1 0 -550 0 1 6600
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_13
timestamp 1675433017
transform 0 -1 7700 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_14
timestamp 1675433017
transform 1 0 -550 0 1 7700
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_15
timestamp 1675433017
transform 0 -1 8800 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_16
timestamp 1675433017
transform 1 0 -550 0 1 8800
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_17
timestamp 1675433017
transform 0 -1 9900 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_18
timestamp 1675433017
transform 1 0 -550 0 1 9900
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_19
timestamp 1675433017
transform 0 -1 11000 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_20
timestamp 1675433017
transform 1 0 -550 0 1 11000
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_21
timestamp 1675433017
transform 0 -1 12100 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_22
timestamp 1675433017
transform 1 0 -550 0 1 12100
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_23
timestamp 1675433017
transform 0 -1 13200 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_24
timestamp 1675433017
transform 1 0 -550 0 1 13200
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_25
timestamp 1675433017
transform 0 -1 14300 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_26
timestamp 1675433017
transform 1 0 -550 0 1 14300
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_27
timestamp 1675433017
transform 0 -1 15400 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_28
timestamp 1675433017
transform 1 0 -550 0 1 15400
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_29
timestamp 1675433017
transform 0 -1 16500 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_30
timestamp 1675433017
transform 1 0 -550 0 1 16500
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_31
timestamp 1675433017
transform 0 -1 17600 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_32
timestamp 1675433017
transform 1 0 -550 0 1 17600
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_33
timestamp 1675433017
transform 0 -1 18700 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_34
timestamp 1675433017
transform 1 0 -550 0 1 18700
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_35
timestamp 1675433017
transform 0 -1 19800 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_36
timestamp 1675433017
transform 1 0 -550 0 1 19800
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_37
timestamp 1675433017
transform 0 -1 20900 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_38
timestamp 1675433017
transform 1 0 -550 0 1 20900
box -975 -113 663 663
use pmos_drain_frame_lt  pmos_drain_frame_lt_39
timestamp 1675433017
transform 0 -1 22000 -1 0 22550
box -975 -113 663 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_0 waffle_cells
timestamp 1675433101
transform 0 -1 550 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_1
timestamp 1675433101
transform 1 0 22000 0 1 550
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_2
timestamp 1675433101
transform 0 -1 1650 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_3
timestamp 1675433101
transform 1 0 22000 0 1 1650
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_4
timestamp 1675433101
transform 0 -1 2750 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_5
timestamp 1675433101
transform 1 0 22000 0 1 2750
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_6
timestamp 1675433101
transform 0 -1 3850 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_7
timestamp 1675433101
transform 1 0 22000 0 1 3850
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_8
timestamp 1675433101
transform 0 -1 4950 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_9
timestamp 1675433101
transform 1 0 22000 0 1 4950
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_10
timestamp 1675433101
transform 0 -1 6050 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_11
timestamp 1675433101
transform 1 0 22000 0 1 6050
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_12
timestamp 1675433101
transform 0 -1 7150 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_13
timestamp 1675433101
transform 1 0 22000 0 1 7150
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_14
timestamp 1675433101
transform 0 -1 8250 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_15
timestamp 1675433101
transform 1 0 22000 0 1 8250
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_16
timestamp 1675433101
transform 0 -1 9350 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_17
timestamp 1675433101
transform 1 0 22000 0 1 9350
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_18
timestamp 1675433101
transform 0 -1 10450 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_19
timestamp 1675433101
transform 1 0 22000 0 1 10450
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_20
timestamp 1675433101
transform 0 -1 11550 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_21
timestamp 1675433101
transform 1 0 22000 0 1 11550
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_22
timestamp 1675433101
transform 0 -1 12650 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_23
timestamp 1675433101
transform 1 0 22000 0 1 12650
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_24
timestamp 1675433101
transform 0 -1 13750 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_25
timestamp 1675433101
transform 1 0 22000 0 1 13750
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_26
timestamp 1675433101
transform 0 -1 14850 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_27
timestamp 1675433101
transform 1 0 22000 0 1 14850
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_28
timestamp 1675433101
transform 0 -1 15950 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_29
timestamp 1675433101
transform 1 0 22000 0 1 15950
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_30
timestamp 1675433101
transform 0 -1 17050 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_31
timestamp 1675433101
transform 1 0 22000 0 1 17050
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_32
timestamp 1675433101
transform 0 -1 18150 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_33
timestamp 1675433101
transform 1 0 22000 0 1 18150
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_34
timestamp 1675433101
transform 0 -1 19250 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_35
timestamp 1675433101
transform 1 0 22000 0 1 19250
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_36
timestamp 1675433101
transform 0 -1 20350 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_37
timestamp 1675433101
transform 1 0 22000 0 1 20350
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_38
timestamp 1675433101
transform 0 -1 21450 -1 0 0
box -113 -113 1575 663
use pmos_drain_frame_rb  pmos_drain_frame_rb_39
timestamp 1675433101
transform 1 0 22000 0 1 21450
box -113 -113 1575 663
use pmos_drain_in  pmos_drain_in_0 waffle_cells
timestamp 1675432984
transform 1 0 0 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_1
timestamp 1675432984
transform 1 0 0 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_2
timestamp 1675432984
transform 1 0 0 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_3
timestamp 1675432984
transform 1 0 0 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_4
timestamp 1675432984
transform 1 0 0 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_5
timestamp 1675432984
transform 1 0 0 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_6
timestamp 1675432984
transform 1 0 0 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_7
timestamp 1675432984
transform 1 0 0 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_8
timestamp 1675432984
transform 1 0 0 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_9
timestamp 1675432984
transform 1 0 0 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_10
timestamp 1675432984
transform 1 0 0 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_11
timestamp 1675432984
transform 1 0 0 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_12
timestamp 1675432984
transform 1 0 0 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_13
timestamp 1675432984
transform 1 0 0 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_14
timestamp 1675432984
transform 1 0 0 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_15
timestamp 1675432984
transform 1 0 0 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_16
timestamp 1675432984
transform 1 0 0 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_17
timestamp 1675432984
transform 1 0 0 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_18
timestamp 1675432984
transform 1 0 0 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_19
timestamp 1675432984
transform 1 0 0 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_20
timestamp 1675432984
transform 1 0 550 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_21
timestamp 1675432984
transform 1 0 550 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_22
timestamp 1675432984
transform 1 0 550 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_23
timestamp 1675432984
transform 1 0 550 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_24
timestamp 1675432984
transform 1 0 550 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_25
timestamp 1675432984
transform 1 0 550 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_26
timestamp 1675432984
transform 1 0 550 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_27
timestamp 1675432984
transform 1 0 550 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_28
timestamp 1675432984
transform 1 0 550 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_29
timestamp 1675432984
transform 1 0 550 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_30
timestamp 1675432984
transform 1 0 550 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_31
timestamp 1675432984
transform 1 0 550 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_32
timestamp 1675432984
transform 1 0 550 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_33
timestamp 1675432984
transform 1 0 550 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_34
timestamp 1675432984
transform 1 0 550 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_35
timestamp 1675432984
transform 1 0 550 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_36
timestamp 1675432984
transform 1 0 550 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_37
timestamp 1675432984
transform 1 0 550 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_38
timestamp 1675432984
transform 1 0 550 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_39
timestamp 1675432984
transform 1 0 550 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_40
timestamp 1675432984
transform 1 0 1100 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_41
timestamp 1675432984
transform 1 0 1100 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_42
timestamp 1675432984
transform 1 0 1100 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_43
timestamp 1675432984
transform 1 0 1100 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_44
timestamp 1675432984
transform 1 0 1100 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_45
timestamp 1675432984
transform 1 0 1100 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_46
timestamp 1675432984
transform 1 0 1100 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_47
timestamp 1675432984
transform 1 0 1100 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_48
timestamp 1675432984
transform 1 0 1100 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_49
timestamp 1675432984
transform 1 0 1100 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_50
timestamp 1675432984
transform 1 0 1100 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_51
timestamp 1675432984
transform 1 0 1100 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_52
timestamp 1675432984
transform 1 0 1100 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_53
timestamp 1675432984
transform 1 0 1100 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_54
timestamp 1675432984
transform 1 0 1100 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_55
timestamp 1675432984
transform 1 0 1100 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_56
timestamp 1675432984
transform 1 0 1100 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_57
timestamp 1675432984
transform 1 0 1100 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_58
timestamp 1675432984
transform 1 0 1100 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_59
timestamp 1675432984
transform 1 0 1100 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_60
timestamp 1675432984
transform 1 0 1650 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_61
timestamp 1675432984
transform 1 0 1650 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_62
timestamp 1675432984
transform 1 0 1650 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_63
timestamp 1675432984
transform 1 0 1650 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_64
timestamp 1675432984
transform 1 0 1650 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_65
timestamp 1675432984
transform 1 0 1650 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_66
timestamp 1675432984
transform 1 0 1650 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_67
timestamp 1675432984
transform 1 0 1650 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_68
timestamp 1675432984
transform 1 0 1650 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_69
timestamp 1675432984
transform 1 0 1650 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_70
timestamp 1675432984
transform 1 0 1650 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_71
timestamp 1675432984
transform 1 0 1650 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_72
timestamp 1675432984
transform 1 0 1650 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_73
timestamp 1675432984
transform 1 0 1650 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_74
timestamp 1675432984
transform 1 0 1650 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_75
timestamp 1675432984
transform 1 0 1650 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_76
timestamp 1675432984
transform 1 0 1650 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_77
timestamp 1675432984
transform 1 0 1650 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_78
timestamp 1675432984
transform 1 0 1650 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_79
timestamp 1675432984
transform 1 0 1650 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_80
timestamp 1675432984
transform 1 0 2200 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_81
timestamp 1675432984
transform 1 0 2200 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_82
timestamp 1675432984
transform 1 0 2200 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_83
timestamp 1675432984
transform 1 0 2200 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_84
timestamp 1675432984
transform 1 0 2200 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_85
timestamp 1675432984
transform 1 0 2200 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_86
timestamp 1675432984
transform 1 0 2200 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_87
timestamp 1675432984
transform 1 0 2200 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_88
timestamp 1675432984
transform 1 0 2200 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_89
timestamp 1675432984
transform 1 0 2200 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_90
timestamp 1675432984
transform 1 0 2200 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_91
timestamp 1675432984
transform 1 0 2200 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_92
timestamp 1675432984
transform 1 0 2200 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_93
timestamp 1675432984
transform 1 0 2200 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_94
timestamp 1675432984
transform 1 0 2200 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_95
timestamp 1675432984
transform 1 0 2200 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_96
timestamp 1675432984
transform 1 0 2200 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_97
timestamp 1675432984
transform 1 0 2200 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_98
timestamp 1675432984
transform 1 0 2200 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_99
timestamp 1675432984
transform 1 0 2200 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_100
timestamp 1675432984
transform 1 0 2750 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_101
timestamp 1675432984
transform 1 0 2750 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_102
timestamp 1675432984
transform 1 0 2750 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_103
timestamp 1675432984
transform 1 0 2750 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_104
timestamp 1675432984
transform 1 0 2750 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_105
timestamp 1675432984
transform 1 0 2750 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_106
timestamp 1675432984
transform 1 0 2750 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_107
timestamp 1675432984
transform 1 0 2750 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_108
timestamp 1675432984
transform 1 0 2750 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_109
timestamp 1675432984
transform 1 0 2750 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_110
timestamp 1675432984
transform 1 0 2750 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_111
timestamp 1675432984
transform 1 0 2750 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_112
timestamp 1675432984
transform 1 0 2750 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_113
timestamp 1675432984
transform 1 0 2750 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_114
timestamp 1675432984
transform 1 0 2750 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_115
timestamp 1675432984
transform 1 0 2750 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_116
timestamp 1675432984
transform 1 0 2750 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_117
timestamp 1675432984
transform 1 0 2750 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_118
timestamp 1675432984
transform 1 0 2750 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_119
timestamp 1675432984
transform 1 0 2750 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_120
timestamp 1675432984
transform 1 0 3300 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_121
timestamp 1675432984
transform 1 0 3300 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_122
timestamp 1675432984
transform 1 0 3300 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_123
timestamp 1675432984
transform 1 0 3300 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_124
timestamp 1675432984
transform 1 0 3300 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_125
timestamp 1675432984
transform 1 0 3300 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_126
timestamp 1675432984
transform 1 0 3300 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_127
timestamp 1675432984
transform 1 0 3300 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_128
timestamp 1675432984
transform 1 0 3300 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_129
timestamp 1675432984
transform 1 0 3300 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_130
timestamp 1675432984
transform 1 0 3300 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_131
timestamp 1675432984
transform 1 0 3300 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_132
timestamp 1675432984
transform 1 0 3300 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_133
timestamp 1675432984
transform 1 0 3300 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_134
timestamp 1675432984
transform 1 0 3300 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_135
timestamp 1675432984
transform 1 0 3300 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_136
timestamp 1675432984
transform 1 0 3300 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_137
timestamp 1675432984
transform 1 0 3300 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_138
timestamp 1675432984
transform 1 0 3300 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_139
timestamp 1675432984
transform 1 0 3300 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_140
timestamp 1675432984
transform 1 0 3850 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_141
timestamp 1675432984
transform 1 0 3850 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_142
timestamp 1675432984
transform 1 0 3850 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_143
timestamp 1675432984
transform 1 0 3850 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_144
timestamp 1675432984
transform 1 0 3850 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_145
timestamp 1675432984
transform 1 0 3850 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_146
timestamp 1675432984
transform 1 0 3850 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_147
timestamp 1675432984
transform 1 0 3850 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_148
timestamp 1675432984
transform 1 0 3850 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_149
timestamp 1675432984
transform 1 0 3850 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_150
timestamp 1675432984
transform 1 0 3850 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_151
timestamp 1675432984
transform 1 0 3850 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_152
timestamp 1675432984
transform 1 0 3850 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_153
timestamp 1675432984
transform 1 0 3850 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_154
timestamp 1675432984
transform 1 0 3850 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_155
timestamp 1675432984
transform 1 0 3850 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_156
timestamp 1675432984
transform 1 0 3850 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_157
timestamp 1675432984
transform 1 0 3850 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_158
timestamp 1675432984
transform 1 0 3850 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_159
timestamp 1675432984
transform 1 0 3850 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_160
timestamp 1675432984
transform 1 0 4400 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_161
timestamp 1675432984
transform 1 0 4400 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_162
timestamp 1675432984
transform 1 0 4400 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_163
timestamp 1675432984
transform 1 0 4400 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_164
timestamp 1675432984
transform 1 0 4400 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_165
timestamp 1675432984
transform 1 0 4400 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_166
timestamp 1675432984
transform 1 0 4400 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_167
timestamp 1675432984
transform 1 0 4400 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_168
timestamp 1675432984
transform 1 0 4400 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_169
timestamp 1675432984
transform 1 0 4400 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_170
timestamp 1675432984
transform 1 0 4400 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_171
timestamp 1675432984
transform 1 0 4400 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_172
timestamp 1675432984
transform 1 0 4400 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_173
timestamp 1675432984
transform 1 0 4400 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_174
timestamp 1675432984
transform 1 0 4400 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_175
timestamp 1675432984
transform 1 0 4400 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_176
timestamp 1675432984
transform 1 0 4400 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_177
timestamp 1675432984
transform 1 0 4400 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_178
timestamp 1675432984
transform 1 0 4400 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_179
timestamp 1675432984
transform 1 0 4400 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_180
timestamp 1675432984
transform 1 0 4950 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_181
timestamp 1675432984
transform 1 0 4950 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_182
timestamp 1675432984
transform 1 0 4950 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_183
timestamp 1675432984
transform 1 0 4950 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_184
timestamp 1675432984
transform 1 0 4950 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_185
timestamp 1675432984
transform 1 0 4950 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_186
timestamp 1675432984
transform 1 0 4950 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_187
timestamp 1675432984
transform 1 0 4950 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_188
timestamp 1675432984
transform 1 0 4950 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_189
timestamp 1675432984
transform 1 0 4950 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_190
timestamp 1675432984
transform 1 0 4950 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_191
timestamp 1675432984
transform 1 0 4950 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_192
timestamp 1675432984
transform 1 0 4950 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_193
timestamp 1675432984
transform 1 0 4950 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_194
timestamp 1675432984
transform 1 0 4950 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_195
timestamp 1675432984
transform 1 0 4950 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_196
timestamp 1675432984
transform 1 0 4950 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_197
timestamp 1675432984
transform 1 0 4950 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_198
timestamp 1675432984
transform 1 0 4950 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_199
timestamp 1675432984
transform 1 0 4950 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_200
timestamp 1675432984
transform 1 0 5500 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_201
timestamp 1675432984
transform 1 0 5500 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_202
timestamp 1675432984
transform 1 0 5500 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_203
timestamp 1675432984
transform 1 0 5500 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_204
timestamp 1675432984
transform 1 0 5500 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_205
timestamp 1675432984
transform 1 0 5500 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_206
timestamp 1675432984
transform 1 0 5500 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_207
timestamp 1675432984
transform 1 0 5500 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_208
timestamp 1675432984
transform 1 0 5500 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_209
timestamp 1675432984
transform 1 0 5500 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_210
timestamp 1675432984
transform 1 0 5500 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_211
timestamp 1675432984
transform 1 0 5500 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_212
timestamp 1675432984
transform 1 0 5500 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_213
timestamp 1675432984
transform 1 0 5500 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_214
timestamp 1675432984
transform 1 0 5500 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_215
timestamp 1675432984
transform 1 0 5500 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_216
timestamp 1675432984
transform 1 0 5500 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_217
timestamp 1675432984
transform 1 0 5500 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_218
timestamp 1675432984
transform 1 0 5500 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_219
timestamp 1675432984
transform 1 0 5500 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_220
timestamp 1675432984
transform 1 0 6050 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_221
timestamp 1675432984
transform 1 0 6050 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_222
timestamp 1675432984
transform 1 0 6050 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_223
timestamp 1675432984
transform 1 0 6050 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_224
timestamp 1675432984
transform 1 0 6050 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_225
timestamp 1675432984
transform 1 0 6050 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_226
timestamp 1675432984
transform 1 0 6050 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_227
timestamp 1675432984
transform 1 0 6050 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_228
timestamp 1675432984
transform 1 0 6050 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_229
timestamp 1675432984
transform 1 0 6050 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_230
timestamp 1675432984
transform 1 0 6050 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_231
timestamp 1675432984
transform 1 0 6050 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_232
timestamp 1675432984
transform 1 0 6050 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_233
timestamp 1675432984
transform 1 0 6050 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_234
timestamp 1675432984
transform 1 0 6050 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_235
timestamp 1675432984
transform 1 0 6050 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_236
timestamp 1675432984
transform 1 0 6050 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_237
timestamp 1675432984
transform 1 0 6050 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_238
timestamp 1675432984
transform 1 0 6050 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_239
timestamp 1675432984
transform 1 0 6050 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_240
timestamp 1675432984
transform 1 0 6600 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_241
timestamp 1675432984
transform 1 0 6600 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_242
timestamp 1675432984
transform 1 0 6600 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_243
timestamp 1675432984
transform 1 0 6600 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_244
timestamp 1675432984
transform 1 0 6600 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_245
timestamp 1675432984
transform 1 0 6600 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_246
timestamp 1675432984
transform 1 0 6600 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_247
timestamp 1675432984
transform 1 0 6600 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_248
timestamp 1675432984
transform 1 0 6600 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_249
timestamp 1675432984
transform 1 0 6600 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_250
timestamp 1675432984
transform 1 0 6600 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_251
timestamp 1675432984
transform 1 0 6600 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_252
timestamp 1675432984
transform 1 0 6600 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_253
timestamp 1675432984
transform 1 0 6600 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_254
timestamp 1675432984
transform 1 0 6600 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_255
timestamp 1675432984
transform 1 0 6600 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_256
timestamp 1675432984
transform 1 0 6600 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_257
timestamp 1675432984
transform 1 0 6600 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_258
timestamp 1675432984
transform 1 0 6600 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_259
timestamp 1675432984
transform 1 0 6600 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_260
timestamp 1675432984
transform 1 0 7150 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_261
timestamp 1675432984
transform 1 0 7150 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_262
timestamp 1675432984
transform 1 0 7150 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_263
timestamp 1675432984
transform 1 0 7150 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_264
timestamp 1675432984
transform 1 0 7150 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_265
timestamp 1675432984
transform 1 0 7150 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_266
timestamp 1675432984
transform 1 0 7150 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_267
timestamp 1675432984
transform 1 0 7150 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_268
timestamp 1675432984
transform 1 0 7150 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_269
timestamp 1675432984
transform 1 0 7150 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_270
timestamp 1675432984
transform 1 0 7150 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_271
timestamp 1675432984
transform 1 0 7150 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_272
timestamp 1675432984
transform 1 0 7150 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_273
timestamp 1675432984
transform 1 0 7150 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_274
timestamp 1675432984
transform 1 0 7150 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_275
timestamp 1675432984
transform 1 0 7150 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_276
timestamp 1675432984
transform 1 0 7150 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_277
timestamp 1675432984
transform 1 0 7150 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_278
timestamp 1675432984
transform 1 0 7150 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_279
timestamp 1675432984
transform 1 0 7150 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_280
timestamp 1675432984
transform 1 0 7700 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_281
timestamp 1675432984
transform 1 0 7700 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_282
timestamp 1675432984
transform 1 0 7700 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_283
timestamp 1675432984
transform 1 0 7700 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_284
timestamp 1675432984
transform 1 0 7700 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_285
timestamp 1675432984
transform 1 0 7700 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_286
timestamp 1675432984
transform 1 0 7700 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_287
timestamp 1675432984
transform 1 0 7700 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_288
timestamp 1675432984
transform 1 0 7700 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_289
timestamp 1675432984
transform 1 0 7700 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_290
timestamp 1675432984
transform 1 0 7700 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_291
timestamp 1675432984
transform 1 0 7700 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_292
timestamp 1675432984
transform 1 0 7700 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_293
timestamp 1675432984
transform 1 0 7700 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_294
timestamp 1675432984
transform 1 0 7700 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_295
timestamp 1675432984
transform 1 0 7700 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_296
timestamp 1675432984
transform 1 0 7700 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_297
timestamp 1675432984
transform 1 0 7700 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_298
timestamp 1675432984
transform 1 0 7700 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_299
timestamp 1675432984
transform 1 0 7700 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_300
timestamp 1675432984
transform 1 0 8250 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_301
timestamp 1675432984
transform 1 0 8250 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_302
timestamp 1675432984
transform 1 0 8250 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_303
timestamp 1675432984
transform 1 0 8250 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_304
timestamp 1675432984
transform 1 0 8250 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_305
timestamp 1675432984
transform 1 0 8250 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_306
timestamp 1675432984
transform 1 0 8250 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_307
timestamp 1675432984
transform 1 0 8250 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_308
timestamp 1675432984
transform 1 0 8250 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_309
timestamp 1675432984
transform 1 0 8250 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_310
timestamp 1675432984
transform 1 0 8250 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_311
timestamp 1675432984
transform 1 0 8250 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_312
timestamp 1675432984
transform 1 0 8250 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_313
timestamp 1675432984
transform 1 0 8250 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_314
timestamp 1675432984
transform 1 0 8250 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_315
timestamp 1675432984
transform 1 0 8250 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_316
timestamp 1675432984
transform 1 0 8250 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_317
timestamp 1675432984
transform 1 0 8250 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_318
timestamp 1675432984
transform 1 0 8250 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_319
timestamp 1675432984
transform 1 0 8250 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_320
timestamp 1675432984
transform 1 0 8800 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_321
timestamp 1675432984
transform 1 0 8800 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_322
timestamp 1675432984
transform 1 0 8800 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_323
timestamp 1675432984
transform 1 0 8800 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_324
timestamp 1675432984
transform 1 0 8800 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_325
timestamp 1675432984
transform 1 0 8800 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_326
timestamp 1675432984
transform 1 0 8800 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_327
timestamp 1675432984
transform 1 0 8800 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_328
timestamp 1675432984
transform 1 0 8800 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_329
timestamp 1675432984
transform 1 0 8800 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_330
timestamp 1675432984
transform 1 0 8800 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_331
timestamp 1675432984
transform 1 0 8800 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_332
timestamp 1675432984
transform 1 0 8800 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_333
timestamp 1675432984
transform 1 0 8800 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_334
timestamp 1675432984
transform 1 0 8800 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_335
timestamp 1675432984
transform 1 0 8800 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_336
timestamp 1675432984
transform 1 0 8800 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_337
timestamp 1675432984
transform 1 0 8800 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_338
timestamp 1675432984
transform 1 0 8800 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_339
timestamp 1675432984
transform 1 0 8800 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_340
timestamp 1675432984
transform 1 0 9350 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_341
timestamp 1675432984
transform 1 0 9350 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_342
timestamp 1675432984
transform 1 0 9350 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_343
timestamp 1675432984
transform 1 0 9350 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_344
timestamp 1675432984
transform 1 0 9350 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_345
timestamp 1675432984
transform 1 0 9350 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_346
timestamp 1675432984
transform 1 0 9350 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_347
timestamp 1675432984
transform 1 0 9350 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_348
timestamp 1675432984
transform 1 0 9350 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_349
timestamp 1675432984
transform 1 0 9350 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_350
timestamp 1675432984
transform 1 0 9350 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_351
timestamp 1675432984
transform 1 0 9350 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_352
timestamp 1675432984
transform 1 0 9350 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_353
timestamp 1675432984
transform 1 0 9350 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_354
timestamp 1675432984
transform 1 0 9350 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_355
timestamp 1675432984
transform 1 0 9350 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_356
timestamp 1675432984
transform 1 0 9350 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_357
timestamp 1675432984
transform 1 0 9350 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_358
timestamp 1675432984
transform 1 0 9350 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_359
timestamp 1675432984
transform 1 0 9350 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_360
timestamp 1675432984
transform 1 0 9900 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_361
timestamp 1675432984
transform 1 0 9900 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_362
timestamp 1675432984
transform 1 0 9900 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_363
timestamp 1675432984
transform 1 0 9900 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_364
timestamp 1675432984
transform 1 0 9900 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_365
timestamp 1675432984
transform 1 0 9900 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_366
timestamp 1675432984
transform 1 0 9900 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_367
timestamp 1675432984
transform 1 0 9900 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_368
timestamp 1675432984
transform 1 0 9900 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_369
timestamp 1675432984
transform 1 0 9900 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_370
timestamp 1675432984
transform 1 0 9900 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_371
timestamp 1675432984
transform 1 0 9900 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_372
timestamp 1675432984
transform 1 0 9900 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_373
timestamp 1675432984
transform 1 0 9900 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_374
timestamp 1675432984
transform 1 0 9900 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_375
timestamp 1675432984
transform 1 0 9900 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_376
timestamp 1675432984
transform 1 0 9900 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_377
timestamp 1675432984
transform 1 0 9900 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_378
timestamp 1675432984
transform 1 0 9900 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_379
timestamp 1675432984
transform 1 0 9900 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_380
timestamp 1675432984
transform 1 0 10450 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_381
timestamp 1675432984
transform 1 0 10450 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_382
timestamp 1675432984
transform 1 0 10450 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_383
timestamp 1675432984
transform 1 0 10450 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_384
timestamp 1675432984
transform 1 0 10450 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_385
timestamp 1675432984
transform 1 0 10450 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_386
timestamp 1675432984
transform 1 0 10450 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_387
timestamp 1675432984
transform 1 0 10450 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_388
timestamp 1675432984
transform 1 0 10450 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_389
timestamp 1675432984
transform 1 0 10450 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_390
timestamp 1675432984
transform 1 0 10450 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_391
timestamp 1675432984
transform 1 0 10450 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_392
timestamp 1675432984
transform 1 0 10450 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_393
timestamp 1675432984
transform 1 0 10450 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_394
timestamp 1675432984
transform 1 0 10450 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_395
timestamp 1675432984
transform 1 0 10450 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_396
timestamp 1675432984
transform 1 0 10450 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_397
timestamp 1675432984
transform 1 0 10450 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_398
timestamp 1675432984
transform 1 0 10450 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_399
timestamp 1675432984
transform 1 0 10450 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_400
timestamp 1675432984
transform 1 0 11000 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_401
timestamp 1675432984
transform 1 0 11000 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_402
timestamp 1675432984
transform 1 0 11000 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_403
timestamp 1675432984
transform 1 0 11000 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_404
timestamp 1675432984
transform 1 0 11000 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_405
timestamp 1675432984
transform 1 0 11000 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_406
timestamp 1675432984
transform 1 0 11000 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_407
timestamp 1675432984
transform 1 0 11000 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_408
timestamp 1675432984
transform 1 0 11000 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_409
timestamp 1675432984
transform 1 0 11000 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_410
timestamp 1675432984
transform 1 0 11000 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_411
timestamp 1675432984
transform 1 0 11000 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_412
timestamp 1675432984
transform 1 0 11000 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_413
timestamp 1675432984
transform 1 0 11000 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_414
timestamp 1675432984
transform 1 0 11000 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_415
timestamp 1675432984
transform 1 0 11000 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_416
timestamp 1675432984
transform 1 0 11000 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_417
timestamp 1675432984
transform 1 0 11000 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_418
timestamp 1675432984
transform 1 0 11000 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_419
timestamp 1675432984
transform 1 0 11000 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_420
timestamp 1675432984
transform 1 0 11550 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_421
timestamp 1675432984
transform 1 0 11550 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_422
timestamp 1675432984
transform 1 0 11550 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_423
timestamp 1675432984
transform 1 0 11550 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_424
timestamp 1675432984
transform 1 0 11550 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_425
timestamp 1675432984
transform 1 0 11550 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_426
timestamp 1675432984
transform 1 0 11550 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_427
timestamp 1675432984
transform 1 0 11550 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_428
timestamp 1675432984
transform 1 0 11550 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_429
timestamp 1675432984
transform 1 0 11550 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_430
timestamp 1675432984
transform 1 0 11550 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_431
timestamp 1675432984
transform 1 0 11550 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_432
timestamp 1675432984
transform 1 0 11550 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_433
timestamp 1675432984
transform 1 0 11550 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_434
timestamp 1675432984
transform 1 0 11550 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_435
timestamp 1675432984
transform 1 0 11550 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_436
timestamp 1675432984
transform 1 0 11550 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_437
timestamp 1675432984
transform 1 0 11550 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_438
timestamp 1675432984
transform 1 0 11550 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_439
timestamp 1675432984
transform 1 0 11550 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_440
timestamp 1675432984
transform 1 0 12100 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_441
timestamp 1675432984
transform 1 0 12100 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_442
timestamp 1675432984
transform 1 0 12100 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_443
timestamp 1675432984
transform 1 0 12100 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_444
timestamp 1675432984
transform 1 0 12100 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_445
timestamp 1675432984
transform 1 0 12100 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_446
timestamp 1675432984
transform 1 0 12100 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_447
timestamp 1675432984
transform 1 0 12100 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_448
timestamp 1675432984
transform 1 0 12100 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_449
timestamp 1675432984
transform 1 0 12100 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_450
timestamp 1675432984
transform 1 0 12100 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_451
timestamp 1675432984
transform 1 0 12100 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_452
timestamp 1675432984
transform 1 0 12100 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_453
timestamp 1675432984
transform 1 0 12100 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_454
timestamp 1675432984
transform 1 0 12100 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_455
timestamp 1675432984
transform 1 0 12100 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_456
timestamp 1675432984
transform 1 0 12100 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_457
timestamp 1675432984
transform 1 0 12100 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_458
timestamp 1675432984
transform 1 0 12100 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_459
timestamp 1675432984
transform 1 0 12100 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_460
timestamp 1675432984
transform 1 0 12650 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_461
timestamp 1675432984
transform 1 0 12650 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_462
timestamp 1675432984
transform 1 0 12650 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_463
timestamp 1675432984
transform 1 0 12650 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_464
timestamp 1675432984
transform 1 0 12650 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_465
timestamp 1675432984
transform 1 0 12650 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_466
timestamp 1675432984
transform 1 0 12650 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_467
timestamp 1675432984
transform 1 0 12650 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_468
timestamp 1675432984
transform 1 0 12650 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_469
timestamp 1675432984
transform 1 0 12650 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_470
timestamp 1675432984
transform 1 0 12650 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_471
timestamp 1675432984
transform 1 0 12650 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_472
timestamp 1675432984
transform 1 0 12650 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_473
timestamp 1675432984
transform 1 0 12650 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_474
timestamp 1675432984
transform 1 0 12650 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_475
timestamp 1675432984
transform 1 0 12650 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_476
timestamp 1675432984
transform 1 0 12650 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_477
timestamp 1675432984
transform 1 0 12650 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_478
timestamp 1675432984
transform 1 0 12650 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_479
timestamp 1675432984
transform 1 0 12650 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_480
timestamp 1675432984
transform 1 0 13200 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_481
timestamp 1675432984
transform 1 0 13200 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_482
timestamp 1675432984
transform 1 0 13200 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_483
timestamp 1675432984
transform 1 0 13200 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_484
timestamp 1675432984
transform 1 0 13200 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_485
timestamp 1675432984
transform 1 0 13200 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_486
timestamp 1675432984
transform 1 0 13200 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_487
timestamp 1675432984
transform 1 0 13200 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_488
timestamp 1675432984
transform 1 0 13200 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_489
timestamp 1675432984
transform 1 0 13200 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_490
timestamp 1675432984
transform 1 0 13200 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_491
timestamp 1675432984
transform 1 0 13200 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_492
timestamp 1675432984
transform 1 0 13200 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_493
timestamp 1675432984
transform 1 0 13200 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_494
timestamp 1675432984
transform 1 0 13200 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_495
timestamp 1675432984
transform 1 0 13200 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_496
timestamp 1675432984
transform 1 0 13200 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_497
timestamp 1675432984
transform 1 0 13200 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_498
timestamp 1675432984
transform 1 0 13200 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_499
timestamp 1675432984
transform 1 0 13200 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_500
timestamp 1675432984
transform 1 0 13750 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_501
timestamp 1675432984
transform 1 0 13750 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_502
timestamp 1675432984
transform 1 0 13750 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_503
timestamp 1675432984
transform 1 0 13750 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_504
timestamp 1675432984
transform 1 0 13750 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_505
timestamp 1675432984
transform 1 0 13750 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_506
timestamp 1675432984
transform 1 0 13750 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_507
timestamp 1675432984
transform 1 0 13750 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_508
timestamp 1675432984
transform 1 0 13750 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_509
timestamp 1675432984
transform 1 0 13750 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_510
timestamp 1675432984
transform 1 0 13750 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_511
timestamp 1675432984
transform 1 0 13750 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_512
timestamp 1675432984
transform 1 0 13750 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_513
timestamp 1675432984
transform 1 0 13750 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_514
timestamp 1675432984
transform 1 0 13750 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_515
timestamp 1675432984
transform 1 0 13750 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_516
timestamp 1675432984
transform 1 0 13750 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_517
timestamp 1675432984
transform 1 0 13750 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_518
timestamp 1675432984
transform 1 0 13750 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_519
timestamp 1675432984
transform 1 0 13750 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_520
timestamp 1675432984
transform 1 0 14300 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_521
timestamp 1675432984
transform 1 0 14300 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_522
timestamp 1675432984
transform 1 0 14300 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_523
timestamp 1675432984
transform 1 0 14300 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_524
timestamp 1675432984
transform 1 0 14300 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_525
timestamp 1675432984
transform 1 0 14300 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_526
timestamp 1675432984
transform 1 0 14300 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_527
timestamp 1675432984
transform 1 0 14300 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_528
timestamp 1675432984
transform 1 0 14300 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_529
timestamp 1675432984
transform 1 0 14300 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_530
timestamp 1675432984
transform 1 0 14300 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_531
timestamp 1675432984
transform 1 0 14300 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_532
timestamp 1675432984
transform 1 0 14300 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_533
timestamp 1675432984
transform 1 0 14300 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_534
timestamp 1675432984
transform 1 0 14300 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_535
timestamp 1675432984
transform 1 0 14300 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_536
timestamp 1675432984
transform 1 0 14300 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_537
timestamp 1675432984
transform 1 0 14300 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_538
timestamp 1675432984
transform 1 0 14300 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_539
timestamp 1675432984
transform 1 0 14300 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_540
timestamp 1675432984
transform 1 0 14850 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_541
timestamp 1675432984
transform 1 0 14850 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_542
timestamp 1675432984
transform 1 0 14850 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_543
timestamp 1675432984
transform 1 0 14850 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_544
timestamp 1675432984
transform 1 0 14850 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_545
timestamp 1675432984
transform 1 0 14850 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_546
timestamp 1675432984
transform 1 0 14850 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_547
timestamp 1675432984
transform 1 0 14850 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_548
timestamp 1675432984
transform 1 0 14850 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_549
timestamp 1675432984
transform 1 0 14850 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_550
timestamp 1675432984
transform 1 0 14850 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_551
timestamp 1675432984
transform 1 0 14850 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_552
timestamp 1675432984
transform 1 0 14850 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_553
timestamp 1675432984
transform 1 0 14850 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_554
timestamp 1675432984
transform 1 0 14850 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_555
timestamp 1675432984
transform 1 0 14850 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_556
timestamp 1675432984
transform 1 0 14850 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_557
timestamp 1675432984
transform 1 0 14850 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_558
timestamp 1675432984
transform 1 0 14850 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_559
timestamp 1675432984
transform 1 0 14850 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_560
timestamp 1675432984
transform 1 0 15400 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_561
timestamp 1675432984
transform 1 0 15400 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_562
timestamp 1675432984
transform 1 0 15400 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_563
timestamp 1675432984
transform 1 0 15400 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_564
timestamp 1675432984
transform 1 0 15400 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_565
timestamp 1675432984
transform 1 0 15400 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_566
timestamp 1675432984
transform 1 0 15400 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_567
timestamp 1675432984
transform 1 0 15400 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_568
timestamp 1675432984
transform 1 0 15400 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_569
timestamp 1675432984
transform 1 0 15400 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_570
timestamp 1675432984
transform 1 0 15400 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_571
timestamp 1675432984
transform 1 0 15400 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_572
timestamp 1675432984
transform 1 0 15400 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_573
timestamp 1675432984
transform 1 0 15400 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_574
timestamp 1675432984
transform 1 0 15400 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_575
timestamp 1675432984
transform 1 0 15400 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_576
timestamp 1675432984
transform 1 0 15400 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_577
timestamp 1675432984
transform 1 0 15400 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_578
timestamp 1675432984
transform 1 0 15400 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_579
timestamp 1675432984
transform 1 0 15400 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_580
timestamp 1675432984
transform 1 0 15950 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_581
timestamp 1675432984
transform 1 0 15950 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_582
timestamp 1675432984
transform 1 0 15950 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_583
timestamp 1675432984
transform 1 0 15950 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_584
timestamp 1675432984
transform 1 0 15950 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_585
timestamp 1675432984
transform 1 0 15950 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_586
timestamp 1675432984
transform 1 0 15950 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_587
timestamp 1675432984
transform 1 0 15950 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_588
timestamp 1675432984
transform 1 0 15950 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_589
timestamp 1675432984
transform 1 0 15950 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_590
timestamp 1675432984
transform 1 0 15950 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_591
timestamp 1675432984
transform 1 0 15950 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_592
timestamp 1675432984
transform 1 0 15950 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_593
timestamp 1675432984
transform 1 0 15950 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_594
timestamp 1675432984
transform 1 0 15950 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_595
timestamp 1675432984
transform 1 0 15950 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_596
timestamp 1675432984
transform 1 0 15950 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_597
timestamp 1675432984
transform 1 0 15950 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_598
timestamp 1675432984
transform 1 0 15950 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_599
timestamp 1675432984
transform 1 0 15950 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_600
timestamp 1675432984
transform 1 0 16500 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_601
timestamp 1675432984
transform 1 0 16500 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_602
timestamp 1675432984
transform 1 0 16500 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_603
timestamp 1675432984
transform 1 0 16500 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_604
timestamp 1675432984
transform 1 0 16500 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_605
timestamp 1675432984
transform 1 0 16500 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_606
timestamp 1675432984
transform 1 0 16500 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_607
timestamp 1675432984
transform 1 0 16500 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_608
timestamp 1675432984
transform 1 0 16500 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_609
timestamp 1675432984
transform 1 0 16500 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_610
timestamp 1675432984
transform 1 0 16500 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_611
timestamp 1675432984
transform 1 0 16500 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_612
timestamp 1675432984
transform 1 0 16500 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_613
timestamp 1675432984
transform 1 0 16500 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_614
timestamp 1675432984
transform 1 0 16500 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_615
timestamp 1675432984
transform 1 0 16500 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_616
timestamp 1675432984
transform 1 0 16500 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_617
timestamp 1675432984
transform 1 0 16500 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_618
timestamp 1675432984
transform 1 0 16500 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_619
timestamp 1675432984
transform 1 0 16500 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_620
timestamp 1675432984
transform 1 0 17050 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_621
timestamp 1675432984
transform 1 0 17050 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_622
timestamp 1675432984
transform 1 0 17050 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_623
timestamp 1675432984
transform 1 0 17050 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_624
timestamp 1675432984
transform 1 0 17050 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_625
timestamp 1675432984
transform 1 0 17050 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_626
timestamp 1675432984
transform 1 0 17050 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_627
timestamp 1675432984
transform 1 0 17050 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_628
timestamp 1675432984
transform 1 0 17050 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_629
timestamp 1675432984
transform 1 0 17050 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_630
timestamp 1675432984
transform 1 0 17050 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_631
timestamp 1675432984
transform 1 0 17050 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_632
timestamp 1675432984
transform 1 0 17050 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_633
timestamp 1675432984
transform 1 0 17050 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_634
timestamp 1675432984
transform 1 0 17050 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_635
timestamp 1675432984
transform 1 0 17050 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_636
timestamp 1675432984
transform 1 0 17050 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_637
timestamp 1675432984
transform 1 0 17050 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_638
timestamp 1675432984
transform 1 0 17050 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_639
timestamp 1675432984
transform 1 0 17050 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_640
timestamp 1675432984
transform 1 0 17600 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_641
timestamp 1675432984
transform 1 0 17600 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_642
timestamp 1675432984
transform 1 0 17600 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_643
timestamp 1675432984
transform 1 0 17600 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_644
timestamp 1675432984
transform 1 0 17600 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_645
timestamp 1675432984
transform 1 0 17600 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_646
timestamp 1675432984
transform 1 0 17600 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_647
timestamp 1675432984
transform 1 0 17600 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_648
timestamp 1675432984
transform 1 0 17600 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_649
timestamp 1675432984
transform 1 0 17600 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_650
timestamp 1675432984
transform 1 0 17600 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_651
timestamp 1675432984
transform 1 0 17600 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_652
timestamp 1675432984
transform 1 0 17600 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_653
timestamp 1675432984
transform 1 0 17600 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_654
timestamp 1675432984
transform 1 0 17600 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_655
timestamp 1675432984
transform 1 0 17600 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_656
timestamp 1675432984
transform 1 0 17600 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_657
timestamp 1675432984
transform 1 0 17600 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_658
timestamp 1675432984
transform 1 0 17600 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_659
timestamp 1675432984
transform 1 0 17600 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_660
timestamp 1675432984
transform 1 0 18150 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_661
timestamp 1675432984
transform 1 0 18150 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_662
timestamp 1675432984
transform 1 0 18150 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_663
timestamp 1675432984
transform 1 0 18150 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_664
timestamp 1675432984
transform 1 0 18150 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_665
timestamp 1675432984
transform 1 0 18150 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_666
timestamp 1675432984
transform 1 0 18150 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_667
timestamp 1675432984
transform 1 0 18150 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_668
timestamp 1675432984
transform 1 0 18150 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_669
timestamp 1675432984
transform 1 0 18150 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_670
timestamp 1675432984
transform 1 0 18150 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_671
timestamp 1675432984
transform 1 0 18150 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_672
timestamp 1675432984
transform 1 0 18150 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_673
timestamp 1675432984
transform 1 0 18150 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_674
timestamp 1675432984
transform 1 0 18150 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_675
timestamp 1675432984
transform 1 0 18150 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_676
timestamp 1675432984
transform 1 0 18150 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_677
timestamp 1675432984
transform 1 0 18150 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_678
timestamp 1675432984
transform 1 0 18150 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_679
timestamp 1675432984
transform 1 0 18150 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_680
timestamp 1675432984
transform 1 0 18700 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_681
timestamp 1675432984
transform 1 0 18700 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_682
timestamp 1675432984
transform 1 0 18700 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_683
timestamp 1675432984
transform 1 0 18700 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_684
timestamp 1675432984
transform 1 0 18700 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_685
timestamp 1675432984
transform 1 0 18700 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_686
timestamp 1675432984
transform 1 0 18700 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_687
timestamp 1675432984
transform 1 0 18700 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_688
timestamp 1675432984
transform 1 0 18700 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_689
timestamp 1675432984
transform 1 0 18700 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_690
timestamp 1675432984
transform 1 0 18700 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_691
timestamp 1675432984
transform 1 0 18700 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_692
timestamp 1675432984
transform 1 0 18700 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_693
timestamp 1675432984
transform 1 0 18700 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_694
timestamp 1675432984
transform 1 0 18700 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_695
timestamp 1675432984
transform 1 0 18700 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_696
timestamp 1675432984
transform 1 0 18700 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_697
timestamp 1675432984
transform 1 0 18700 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_698
timestamp 1675432984
transform 1 0 18700 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_699
timestamp 1675432984
transform 1 0 18700 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_700
timestamp 1675432984
transform 1 0 19250 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_701
timestamp 1675432984
transform 1 0 19250 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_702
timestamp 1675432984
transform 1 0 19250 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_703
timestamp 1675432984
transform 1 0 19250 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_704
timestamp 1675432984
transform 1 0 19250 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_705
timestamp 1675432984
transform 1 0 19250 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_706
timestamp 1675432984
transform 1 0 19250 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_707
timestamp 1675432984
transform 1 0 19250 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_708
timestamp 1675432984
transform 1 0 19250 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_709
timestamp 1675432984
transform 1 0 19250 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_710
timestamp 1675432984
transform 1 0 19250 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_711
timestamp 1675432984
transform 1 0 19250 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_712
timestamp 1675432984
transform 1 0 19250 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_713
timestamp 1675432984
transform 1 0 19250 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_714
timestamp 1675432984
transform 1 0 19250 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_715
timestamp 1675432984
transform 1 0 19250 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_716
timestamp 1675432984
transform 1 0 19250 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_717
timestamp 1675432984
transform 1 0 19250 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_718
timestamp 1675432984
transform 1 0 19250 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_719
timestamp 1675432984
transform 1 0 19250 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_720
timestamp 1675432984
transform 1 0 19800 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_721
timestamp 1675432984
transform 1 0 19800 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_722
timestamp 1675432984
transform 1 0 19800 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_723
timestamp 1675432984
transform 1 0 19800 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_724
timestamp 1675432984
transform 1 0 19800 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_725
timestamp 1675432984
transform 1 0 19800 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_726
timestamp 1675432984
transform 1 0 19800 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_727
timestamp 1675432984
transform 1 0 19800 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_728
timestamp 1675432984
transform 1 0 19800 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_729
timestamp 1675432984
transform 1 0 19800 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_730
timestamp 1675432984
transform 1 0 19800 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_731
timestamp 1675432984
transform 1 0 19800 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_732
timestamp 1675432984
transform 1 0 19800 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_733
timestamp 1675432984
transform 1 0 19800 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_734
timestamp 1675432984
transform 1 0 19800 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_735
timestamp 1675432984
transform 1 0 19800 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_736
timestamp 1675432984
transform 1 0 19800 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_737
timestamp 1675432984
transform 1 0 19800 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_738
timestamp 1675432984
transform 1 0 19800 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_739
timestamp 1675432984
transform 1 0 19800 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_740
timestamp 1675432984
transform 1 0 20350 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_741
timestamp 1675432984
transform 1 0 20350 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_742
timestamp 1675432984
transform 1 0 20350 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_743
timestamp 1675432984
transform 1 0 20350 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_744
timestamp 1675432984
transform 1 0 20350 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_745
timestamp 1675432984
transform 1 0 20350 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_746
timestamp 1675432984
transform 1 0 20350 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_747
timestamp 1675432984
transform 1 0 20350 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_748
timestamp 1675432984
transform 1 0 20350 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_749
timestamp 1675432984
transform 1 0 20350 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_750
timestamp 1675432984
transform 1 0 20350 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_751
timestamp 1675432984
transform 1 0 20350 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_752
timestamp 1675432984
transform 1 0 20350 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_753
timestamp 1675432984
transform 1 0 20350 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_754
timestamp 1675432984
transform 1 0 20350 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_755
timestamp 1675432984
transform 1 0 20350 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_756
timestamp 1675432984
transform 1 0 20350 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_757
timestamp 1675432984
transform 1 0 20350 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_758
timestamp 1675432984
transform 1 0 20350 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_759
timestamp 1675432984
transform 1 0 20350 0 1 20900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_760
timestamp 1675432984
transform 1 0 20900 0 1 550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_761
timestamp 1675432984
transform 1 0 20900 0 1 1650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_762
timestamp 1675432984
transform 1 0 20900 0 1 2750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_763
timestamp 1675432984
transform 1 0 20900 0 1 3850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_764
timestamp 1675432984
transform 1 0 20900 0 1 4950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_765
timestamp 1675432984
transform 1 0 20900 0 1 6050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_766
timestamp 1675432984
transform 1 0 20900 0 1 7150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_767
timestamp 1675432984
transform 1 0 20900 0 1 8250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_768
timestamp 1675432984
transform 1 0 20900 0 1 9350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_769
timestamp 1675432984
transform 1 0 20900 0 1 10450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_770
timestamp 1675432984
transform 1 0 20900 0 1 11550
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_771
timestamp 1675432984
transform 1 0 20900 0 1 12650
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_772
timestamp 1675432984
transform 1 0 20900 0 1 13750
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_773
timestamp 1675432984
transform 1 0 20900 0 1 14850
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_774
timestamp 1675432984
transform 1 0 20900 0 1 15950
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_775
timestamp 1675432984
transform 1 0 20900 0 1 17050
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_776
timestamp 1675432984
transform 1 0 20900 0 1 18150
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_777
timestamp 1675432984
transform 1 0 20900 0 1 19250
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_778
timestamp 1675432984
transform 1 0 20900 0 1 20350
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_779
timestamp 1675432984
transform 1 0 20900 0 1 21450
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_780
timestamp 1675432984
transform 1 0 21450 0 1 0
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_781
timestamp 1675432984
transform 1 0 21450 0 1 1100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_782
timestamp 1675432984
transform 1 0 21450 0 1 2200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_783
timestamp 1675432984
transform 1 0 21450 0 1 3300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_784
timestamp 1675432984
transform 1 0 21450 0 1 4400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_785
timestamp 1675432984
transform 1 0 21450 0 1 5500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_786
timestamp 1675432984
transform 1 0 21450 0 1 6600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_787
timestamp 1675432984
transform 1 0 21450 0 1 7700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_788
timestamp 1675432984
transform 1 0 21450 0 1 8800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_789
timestamp 1675432984
transform 1 0 21450 0 1 9900
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_790
timestamp 1675432984
transform 1 0 21450 0 1 11000
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_791
timestamp 1675432984
transform 1 0 21450 0 1 12100
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_792
timestamp 1675432984
transform 1 0 21450 0 1 13200
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_793
timestamp 1675432984
transform 1 0 21450 0 1 14300
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_794
timestamp 1675432984
transform 1 0 21450 0 1 15400
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_795
timestamp 1675432984
transform 1 0 21450 0 1 16500
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_796
timestamp 1675432984
transform 1 0 21450 0 1 17600
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_797
timestamp 1675432984
transform 1 0 21450 0 1 18700
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_798
timestamp 1675432984
transform 1 0 21450 0 1 19800
box -113 -113 663 663
use pmos_drain_in  pmos_drain_in_799
timestamp 1675432984
transform 1 0 21450 0 1 20900
box -113 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_0 waffle_cells
timestamp 1675433049
transform 0 -1 550 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_1
timestamp 1675433049
transform 1 0 -550 0 1 550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_2
timestamp 1675433049
transform 0 -1 1650 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_3
timestamp 1675433049
transform 1 0 -550 0 1 1650
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_4
timestamp 1675433049
transform 0 -1 2750 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_5
timestamp 1675433049
transform 1 0 -550 0 1 2750
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_6
timestamp 1675433049
transform 0 -1 3850 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_7
timestamp 1675433049
transform 1 0 -550 0 1 3850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_8
timestamp 1675433049
transform 0 -1 4950 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_9
timestamp 1675433049
transform 1 0 -550 0 1 4950
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_10
timestamp 1675433049
transform 0 -1 6050 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_11
timestamp 1675433049
transform 1 0 -550 0 1 6050
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_12
timestamp 1675433049
transform 0 -1 7150 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_13
timestamp 1675433049
transform 1 0 -550 0 1 7150
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_14
timestamp 1675433049
transform 0 -1 8250 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_15
timestamp 1675433049
transform 1 0 -550 0 1 8250
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_16
timestamp 1675433049
transform 0 -1 9350 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_17
timestamp 1675433049
transform 1 0 -550 0 1 9350
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_18
timestamp 1675433049
transform 0 -1 10450 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_19
timestamp 1675433049
transform 1 0 -550 0 1 10450
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_20
timestamp 1675433049
transform 0 -1 11550 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_21
timestamp 1675433049
transform 1 0 -550 0 1 11550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_22
timestamp 1675433049
transform 0 -1 12650 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_23
timestamp 1675433049
transform 1 0 -550 0 1 12650
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_24
timestamp 1675433049
transform 0 -1 13750 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_25
timestamp 1675433049
transform 1 0 -550 0 1 13750
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_26
timestamp 1675433049
transform 0 -1 14850 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_27
timestamp 1675433049
transform 1 0 -550 0 1 14850
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_28
timestamp 1675433049
transform 0 -1 15950 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_29
timestamp 1675433049
transform 1 0 -550 0 1 15950
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_30
timestamp 1675433049
transform 0 -1 17050 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_31
timestamp 1675433049
transform 1 0 -550 0 1 17050
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_32
timestamp 1675433049
transform 0 -1 18150 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_33
timestamp 1675433049
transform 1 0 -550 0 1 18150
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_34
timestamp 1675433049
transform 0 -1 19250 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_35
timestamp 1675433049
transform 1 0 -550 0 1 19250
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_36
timestamp 1675433049
transform 0 -1 20350 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_37
timestamp 1675433049
transform 1 0 -550 0 1 20350
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_38
timestamp 1675433049
transform 0 -1 21450 -1 0 22550
box -975 -113 663 663
use pmos_source_frame_lt  pmos_source_frame_lt_39
timestamp 1675433049
transform 1 0 -550 0 1 21450
box -975 -113 663 663
use pmos_source_frame_rb  pmos_source_frame_rb_0 waffle_cells
timestamp 1675433193
transform 1 0 22000 0 1 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_1
timestamp 1675433193
transform 0 -1 1100 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_2
timestamp 1675433193
transform 1 0 22000 0 1 1100
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_3
timestamp 1675433193
transform 0 -1 2200 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_4
timestamp 1675433193
transform 1 0 22000 0 1 2200
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_5
timestamp 1675433193
transform 0 -1 3300 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_6
timestamp 1675433193
transform 1 0 22000 0 1 3300
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_7
timestamp 1675433193
transform 0 -1 4400 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_8
timestamp 1675433193
transform 1 0 22000 0 1 4400
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_9
timestamp 1675433193
transform 0 -1 5500 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_10
timestamp 1675433193
transform 1 0 22000 0 1 5500
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_11
timestamp 1675433193
transform 0 -1 6600 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_12
timestamp 1675433193
transform 1 0 22000 0 1 6600
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_13
timestamp 1675433193
transform 0 -1 7700 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_14
timestamp 1675433193
transform 1 0 22000 0 1 7700
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_15
timestamp 1675433193
transform 0 -1 8800 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_16
timestamp 1675433193
transform 1 0 22000 0 1 8800
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_17
timestamp 1675433193
transform 0 -1 9900 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_18
timestamp 1675433193
transform 1 0 22000 0 1 9900
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_19
timestamp 1675433193
transform 0 -1 11000 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_20
timestamp 1675433193
transform 1 0 22000 0 1 11000
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_21
timestamp 1675433193
transform 0 -1 12100 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_22
timestamp 1675433193
transform 1 0 22000 0 1 12100
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_23
timestamp 1675433193
transform 0 -1 13200 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_24
timestamp 1675433193
transform 1 0 22000 0 1 13200
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_25
timestamp 1675433193
transform 0 -1 14300 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_26
timestamp 1675433193
transform 1 0 22000 0 1 14300
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_27
timestamp 1675433193
transform 0 -1 15400 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_28
timestamp 1675433193
transform 1 0 22000 0 1 15400
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_29
timestamp 1675433193
transform 0 -1 16500 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_30
timestamp 1675433193
transform 1 0 22000 0 1 16500
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_31
timestamp 1675433193
transform 0 -1 17600 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_32
timestamp 1675433193
transform 1 0 22000 0 1 17600
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_33
timestamp 1675433193
transform 0 -1 18700 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_34
timestamp 1675433193
transform 1 0 22000 0 1 18700
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_35
timestamp 1675433193
transform 0 -1 19800 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_36
timestamp 1675433193
transform 1 0 22000 0 1 19800
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_37
timestamp 1675433193
transform 0 -1 20900 -1 0 0
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_38
timestamp 1675433193
transform 1 0 22000 0 1 20900
box -113 -113 1575 663
use pmos_source_frame_rb  pmos_source_frame_rb_39
timestamp 1675433193
transform 0 -1 22000 -1 0 0
box -113 -113 1575 663
use pmos_source_in  pmos_source_in_0 waffle_cells
timestamp 1675432918
transform 1 0 0 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_1
timestamp 1675432918
transform 1 0 0 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_2
timestamp 1675432918
transform 1 0 0 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_3
timestamp 1675432918
transform 1 0 0 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_4
timestamp 1675432918
transform 1 0 0 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_5
timestamp 1675432918
transform 1 0 0 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_6
timestamp 1675432918
transform 1 0 0 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_7
timestamp 1675432918
transform 1 0 0 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_8
timestamp 1675432918
transform 1 0 0 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_9
timestamp 1675432918
transform 1 0 0 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_10
timestamp 1675432918
transform 1 0 0 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_11
timestamp 1675432918
transform 1 0 0 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_12
timestamp 1675432918
transform 1 0 0 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_13
timestamp 1675432918
transform 1 0 0 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_14
timestamp 1675432918
transform 1 0 0 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_15
timestamp 1675432918
transform 1 0 0 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_16
timestamp 1675432918
transform 1 0 0 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_17
timestamp 1675432918
transform 1 0 0 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_18
timestamp 1675432918
transform 1 0 0 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_19
timestamp 1675432918
transform 1 0 0 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_20
timestamp 1675432918
transform 1 0 550 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_21
timestamp 1675432918
transform 1 0 550 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_22
timestamp 1675432918
transform 1 0 550 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_23
timestamp 1675432918
transform 1 0 550 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_24
timestamp 1675432918
transform 1 0 550 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_25
timestamp 1675432918
transform 1 0 550 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_26
timestamp 1675432918
transform 1 0 550 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_27
timestamp 1675432918
transform 1 0 550 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_28
timestamp 1675432918
transform 1 0 550 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_29
timestamp 1675432918
transform 1 0 550 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_30
timestamp 1675432918
transform 1 0 550 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_31
timestamp 1675432918
transform 1 0 550 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_32
timestamp 1675432918
transform 1 0 550 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_33
timestamp 1675432918
transform 1 0 550 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_34
timestamp 1675432918
transform 1 0 550 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_35
timestamp 1675432918
transform 1 0 550 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_36
timestamp 1675432918
transform 1 0 550 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_37
timestamp 1675432918
transform 1 0 550 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_38
timestamp 1675432918
transform 1 0 550 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_39
timestamp 1675432918
transform 1 0 550 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_40
timestamp 1675432918
transform 1 0 1100 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_41
timestamp 1675432918
transform 1 0 1100 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_42
timestamp 1675432918
transform 1 0 1100 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_43
timestamp 1675432918
transform 1 0 1100 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_44
timestamp 1675432918
transform 1 0 1100 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_45
timestamp 1675432918
transform 1 0 1100 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_46
timestamp 1675432918
transform 1 0 1100 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_47
timestamp 1675432918
transform 1 0 1100 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_48
timestamp 1675432918
transform 1 0 1100 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_49
timestamp 1675432918
transform 1 0 1100 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_50
timestamp 1675432918
transform 1 0 1100 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_51
timestamp 1675432918
transform 1 0 1100 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_52
timestamp 1675432918
transform 1 0 1100 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_53
timestamp 1675432918
transform 1 0 1100 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_54
timestamp 1675432918
transform 1 0 1100 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_55
timestamp 1675432918
transform 1 0 1100 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_56
timestamp 1675432918
transform 1 0 1100 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_57
timestamp 1675432918
transform 1 0 1100 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_58
timestamp 1675432918
transform 1 0 1100 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_59
timestamp 1675432918
transform 1 0 1100 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_60
timestamp 1675432918
transform 1 0 1650 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_61
timestamp 1675432918
transform 1 0 1650 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_62
timestamp 1675432918
transform 1 0 1650 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_63
timestamp 1675432918
transform 1 0 1650 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_64
timestamp 1675432918
transform 1 0 1650 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_65
timestamp 1675432918
transform 1 0 1650 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_66
timestamp 1675432918
transform 1 0 1650 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_67
timestamp 1675432918
transform 1 0 1650 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_68
timestamp 1675432918
transform 1 0 1650 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_69
timestamp 1675432918
transform 1 0 1650 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_70
timestamp 1675432918
transform 1 0 1650 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_71
timestamp 1675432918
transform 1 0 1650 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_72
timestamp 1675432918
transform 1 0 1650 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_73
timestamp 1675432918
transform 1 0 1650 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_74
timestamp 1675432918
transform 1 0 1650 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_75
timestamp 1675432918
transform 1 0 1650 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_76
timestamp 1675432918
transform 1 0 1650 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_77
timestamp 1675432918
transform 1 0 1650 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_78
timestamp 1675432918
transform 1 0 1650 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_79
timestamp 1675432918
transform 1 0 1650 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_80
timestamp 1675432918
transform 1 0 2200 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_81
timestamp 1675432918
transform 1 0 2200 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_82
timestamp 1675432918
transform 1 0 2200 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_83
timestamp 1675432918
transform 1 0 2200 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_84
timestamp 1675432918
transform 1 0 2200 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_85
timestamp 1675432918
transform 1 0 2200 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_86
timestamp 1675432918
transform 1 0 2200 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_87
timestamp 1675432918
transform 1 0 2200 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_88
timestamp 1675432918
transform 1 0 2200 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_89
timestamp 1675432918
transform 1 0 2200 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_90
timestamp 1675432918
transform 1 0 2200 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_91
timestamp 1675432918
transform 1 0 2200 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_92
timestamp 1675432918
transform 1 0 2200 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_93
timestamp 1675432918
transform 1 0 2200 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_94
timestamp 1675432918
transform 1 0 2200 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_95
timestamp 1675432918
transform 1 0 2200 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_96
timestamp 1675432918
transform 1 0 2200 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_97
timestamp 1675432918
transform 1 0 2200 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_98
timestamp 1675432918
transform 1 0 2200 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_99
timestamp 1675432918
transform 1 0 2200 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_100
timestamp 1675432918
transform 1 0 2750 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_101
timestamp 1675432918
transform 1 0 2750 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_102
timestamp 1675432918
transform 1 0 2750 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_103
timestamp 1675432918
transform 1 0 2750 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_104
timestamp 1675432918
transform 1 0 2750 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_105
timestamp 1675432918
transform 1 0 2750 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_106
timestamp 1675432918
transform 1 0 2750 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_107
timestamp 1675432918
transform 1 0 2750 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_108
timestamp 1675432918
transform 1 0 2750 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_109
timestamp 1675432918
transform 1 0 2750 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_110
timestamp 1675432918
transform 1 0 2750 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_111
timestamp 1675432918
transform 1 0 2750 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_112
timestamp 1675432918
transform 1 0 2750 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_113
timestamp 1675432918
transform 1 0 2750 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_114
timestamp 1675432918
transform 1 0 2750 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_115
timestamp 1675432918
transform 1 0 2750 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_116
timestamp 1675432918
transform 1 0 2750 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_117
timestamp 1675432918
transform 1 0 2750 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_118
timestamp 1675432918
transform 1 0 2750 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_119
timestamp 1675432918
transform 1 0 2750 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_120
timestamp 1675432918
transform 1 0 3300 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_121
timestamp 1675432918
transform 1 0 3300 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_122
timestamp 1675432918
transform 1 0 3300 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_123
timestamp 1675432918
transform 1 0 3300 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_124
timestamp 1675432918
transform 1 0 3300 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_125
timestamp 1675432918
transform 1 0 3300 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_126
timestamp 1675432918
transform 1 0 3300 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_127
timestamp 1675432918
transform 1 0 3300 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_128
timestamp 1675432918
transform 1 0 3300 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_129
timestamp 1675432918
transform 1 0 3300 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_130
timestamp 1675432918
transform 1 0 3300 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_131
timestamp 1675432918
transform 1 0 3300 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_132
timestamp 1675432918
transform 1 0 3300 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_133
timestamp 1675432918
transform 1 0 3300 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_134
timestamp 1675432918
transform 1 0 3300 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_135
timestamp 1675432918
transform 1 0 3300 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_136
timestamp 1675432918
transform 1 0 3300 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_137
timestamp 1675432918
transform 1 0 3300 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_138
timestamp 1675432918
transform 1 0 3300 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_139
timestamp 1675432918
transform 1 0 3300 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_140
timestamp 1675432918
transform 1 0 3850 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_141
timestamp 1675432918
transform 1 0 3850 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_142
timestamp 1675432918
transform 1 0 3850 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_143
timestamp 1675432918
transform 1 0 3850 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_144
timestamp 1675432918
transform 1 0 3850 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_145
timestamp 1675432918
transform 1 0 3850 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_146
timestamp 1675432918
transform 1 0 3850 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_147
timestamp 1675432918
transform 1 0 3850 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_148
timestamp 1675432918
transform 1 0 3850 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_149
timestamp 1675432918
transform 1 0 3850 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_150
timestamp 1675432918
transform 1 0 3850 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_151
timestamp 1675432918
transform 1 0 3850 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_152
timestamp 1675432918
transform 1 0 3850 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_153
timestamp 1675432918
transform 1 0 3850 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_154
timestamp 1675432918
transform 1 0 3850 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_155
timestamp 1675432918
transform 1 0 3850 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_156
timestamp 1675432918
transform 1 0 3850 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_157
timestamp 1675432918
transform 1 0 3850 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_158
timestamp 1675432918
transform 1 0 3850 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_159
timestamp 1675432918
transform 1 0 3850 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_160
timestamp 1675432918
transform 1 0 4400 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_161
timestamp 1675432918
transform 1 0 4400 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_162
timestamp 1675432918
transform 1 0 4400 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_163
timestamp 1675432918
transform 1 0 4400 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_164
timestamp 1675432918
transform 1 0 4400 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_165
timestamp 1675432918
transform 1 0 4400 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_166
timestamp 1675432918
transform 1 0 4400 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_167
timestamp 1675432918
transform 1 0 4400 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_168
timestamp 1675432918
transform 1 0 4400 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_169
timestamp 1675432918
transform 1 0 4400 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_170
timestamp 1675432918
transform 1 0 4400 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_171
timestamp 1675432918
transform 1 0 4400 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_172
timestamp 1675432918
transform 1 0 4400 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_173
timestamp 1675432918
transform 1 0 4400 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_174
timestamp 1675432918
transform 1 0 4400 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_175
timestamp 1675432918
transform 1 0 4400 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_176
timestamp 1675432918
transform 1 0 4400 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_177
timestamp 1675432918
transform 1 0 4400 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_178
timestamp 1675432918
transform 1 0 4400 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_179
timestamp 1675432918
transform 1 0 4400 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_180
timestamp 1675432918
transform 1 0 4950 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_181
timestamp 1675432918
transform 1 0 4950 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_182
timestamp 1675432918
transform 1 0 4950 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_183
timestamp 1675432918
transform 1 0 4950 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_184
timestamp 1675432918
transform 1 0 4950 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_185
timestamp 1675432918
transform 1 0 4950 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_186
timestamp 1675432918
transform 1 0 4950 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_187
timestamp 1675432918
transform 1 0 4950 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_188
timestamp 1675432918
transform 1 0 4950 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_189
timestamp 1675432918
transform 1 0 4950 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_190
timestamp 1675432918
transform 1 0 4950 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_191
timestamp 1675432918
transform 1 0 4950 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_192
timestamp 1675432918
transform 1 0 4950 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_193
timestamp 1675432918
transform 1 0 4950 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_194
timestamp 1675432918
transform 1 0 4950 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_195
timestamp 1675432918
transform 1 0 4950 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_196
timestamp 1675432918
transform 1 0 4950 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_197
timestamp 1675432918
transform 1 0 4950 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_198
timestamp 1675432918
transform 1 0 4950 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_199
timestamp 1675432918
transform 1 0 4950 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_200
timestamp 1675432918
transform 1 0 5500 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_201
timestamp 1675432918
transform 1 0 5500 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_202
timestamp 1675432918
transform 1 0 5500 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_203
timestamp 1675432918
transform 1 0 5500 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_204
timestamp 1675432918
transform 1 0 5500 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_205
timestamp 1675432918
transform 1 0 5500 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_206
timestamp 1675432918
transform 1 0 5500 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_207
timestamp 1675432918
transform 1 0 5500 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_208
timestamp 1675432918
transform 1 0 5500 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_209
timestamp 1675432918
transform 1 0 5500 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_210
timestamp 1675432918
transform 1 0 5500 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_211
timestamp 1675432918
transform 1 0 5500 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_212
timestamp 1675432918
transform 1 0 5500 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_213
timestamp 1675432918
transform 1 0 5500 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_214
timestamp 1675432918
transform 1 0 5500 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_215
timestamp 1675432918
transform 1 0 5500 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_216
timestamp 1675432918
transform 1 0 5500 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_217
timestamp 1675432918
transform 1 0 5500 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_218
timestamp 1675432918
transform 1 0 5500 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_219
timestamp 1675432918
transform 1 0 5500 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_220
timestamp 1675432918
transform 1 0 6050 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_221
timestamp 1675432918
transform 1 0 6050 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_222
timestamp 1675432918
transform 1 0 6050 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_223
timestamp 1675432918
transform 1 0 6050 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_224
timestamp 1675432918
transform 1 0 6050 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_225
timestamp 1675432918
transform 1 0 6050 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_226
timestamp 1675432918
transform 1 0 6050 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_227
timestamp 1675432918
transform 1 0 6050 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_228
timestamp 1675432918
transform 1 0 6050 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_229
timestamp 1675432918
transform 1 0 6050 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_230
timestamp 1675432918
transform 1 0 6050 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_231
timestamp 1675432918
transform 1 0 6050 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_232
timestamp 1675432918
transform 1 0 6050 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_233
timestamp 1675432918
transform 1 0 6050 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_234
timestamp 1675432918
transform 1 0 6050 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_235
timestamp 1675432918
transform 1 0 6050 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_236
timestamp 1675432918
transform 1 0 6050 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_237
timestamp 1675432918
transform 1 0 6050 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_238
timestamp 1675432918
transform 1 0 6050 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_239
timestamp 1675432918
transform 1 0 6050 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_240
timestamp 1675432918
transform 1 0 6600 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_241
timestamp 1675432918
transform 1 0 6600 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_242
timestamp 1675432918
transform 1 0 6600 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_243
timestamp 1675432918
transform 1 0 6600 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_244
timestamp 1675432918
transform 1 0 6600 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_245
timestamp 1675432918
transform 1 0 6600 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_246
timestamp 1675432918
transform 1 0 6600 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_247
timestamp 1675432918
transform 1 0 6600 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_248
timestamp 1675432918
transform 1 0 6600 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_249
timestamp 1675432918
transform 1 0 6600 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_250
timestamp 1675432918
transform 1 0 6600 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_251
timestamp 1675432918
transform 1 0 6600 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_252
timestamp 1675432918
transform 1 0 6600 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_253
timestamp 1675432918
transform 1 0 6600 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_254
timestamp 1675432918
transform 1 0 6600 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_255
timestamp 1675432918
transform 1 0 6600 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_256
timestamp 1675432918
transform 1 0 6600 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_257
timestamp 1675432918
transform 1 0 6600 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_258
timestamp 1675432918
transform 1 0 6600 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_259
timestamp 1675432918
transform 1 0 6600 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_260
timestamp 1675432918
transform 1 0 7150 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_261
timestamp 1675432918
transform 1 0 7150 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_262
timestamp 1675432918
transform 1 0 7150 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_263
timestamp 1675432918
transform 1 0 7150 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_264
timestamp 1675432918
transform 1 0 7150 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_265
timestamp 1675432918
transform 1 0 7150 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_266
timestamp 1675432918
transform 1 0 7150 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_267
timestamp 1675432918
transform 1 0 7150 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_268
timestamp 1675432918
transform 1 0 7150 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_269
timestamp 1675432918
transform 1 0 7150 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_270
timestamp 1675432918
transform 1 0 7150 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_271
timestamp 1675432918
transform 1 0 7150 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_272
timestamp 1675432918
transform 1 0 7150 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_273
timestamp 1675432918
transform 1 0 7150 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_274
timestamp 1675432918
transform 1 0 7150 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_275
timestamp 1675432918
transform 1 0 7150 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_276
timestamp 1675432918
transform 1 0 7150 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_277
timestamp 1675432918
transform 1 0 7150 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_278
timestamp 1675432918
transform 1 0 7150 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_279
timestamp 1675432918
transform 1 0 7150 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_280
timestamp 1675432918
transform 1 0 7700 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_281
timestamp 1675432918
transform 1 0 7700 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_282
timestamp 1675432918
transform 1 0 7700 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_283
timestamp 1675432918
transform 1 0 7700 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_284
timestamp 1675432918
transform 1 0 7700 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_285
timestamp 1675432918
transform 1 0 7700 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_286
timestamp 1675432918
transform 1 0 7700 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_287
timestamp 1675432918
transform 1 0 7700 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_288
timestamp 1675432918
transform 1 0 7700 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_289
timestamp 1675432918
transform 1 0 7700 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_290
timestamp 1675432918
transform 1 0 7700 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_291
timestamp 1675432918
transform 1 0 7700 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_292
timestamp 1675432918
transform 1 0 7700 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_293
timestamp 1675432918
transform 1 0 7700 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_294
timestamp 1675432918
transform 1 0 7700 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_295
timestamp 1675432918
transform 1 0 7700 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_296
timestamp 1675432918
transform 1 0 7700 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_297
timestamp 1675432918
transform 1 0 7700 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_298
timestamp 1675432918
transform 1 0 7700 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_299
timestamp 1675432918
transform 1 0 7700 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_300
timestamp 1675432918
transform 1 0 8250 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_301
timestamp 1675432918
transform 1 0 8250 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_302
timestamp 1675432918
transform 1 0 8250 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_303
timestamp 1675432918
transform 1 0 8250 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_304
timestamp 1675432918
transform 1 0 8250 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_305
timestamp 1675432918
transform 1 0 8250 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_306
timestamp 1675432918
transform 1 0 8250 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_307
timestamp 1675432918
transform 1 0 8250 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_308
timestamp 1675432918
transform 1 0 8250 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_309
timestamp 1675432918
transform 1 0 8250 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_310
timestamp 1675432918
transform 1 0 8250 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_311
timestamp 1675432918
transform 1 0 8250 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_312
timestamp 1675432918
transform 1 0 8250 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_313
timestamp 1675432918
transform 1 0 8250 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_314
timestamp 1675432918
transform 1 0 8250 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_315
timestamp 1675432918
transform 1 0 8250 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_316
timestamp 1675432918
transform 1 0 8250 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_317
timestamp 1675432918
transform 1 0 8250 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_318
timestamp 1675432918
transform 1 0 8250 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_319
timestamp 1675432918
transform 1 0 8250 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_320
timestamp 1675432918
transform 1 0 8800 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_321
timestamp 1675432918
transform 1 0 8800 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_322
timestamp 1675432918
transform 1 0 8800 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_323
timestamp 1675432918
transform 1 0 8800 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_324
timestamp 1675432918
transform 1 0 8800 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_325
timestamp 1675432918
transform 1 0 8800 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_326
timestamp 1675432918
transform 1 0 8800 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_327
timestamp 1675432918
transform 1 0 8800 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_328
timestamp 1675432918
transform 1 0 8800 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_329
timestamp 1675432918
transform 1 0 8800 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_330
timestamp 1675432918
transform 1 0 8800 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_331
timestamp 1675432918
transform 1 0 8800 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_332
timestamp 1675432918
transform 1 0 8800 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_333
timestamp 1675432918
transform 1 0 8800 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_334
timestamp 1675432918
transform 1 0 8800 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_335
timestamp 1675432918
transform 1 0 8800 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_336
timestamp 1675432918
transform 1 0 8800 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_337
timestamp 1675432918
transform 1 0 8800 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_338
timestamp 1675432918
transform 1 0 8800 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_339
timestamp 1675432918
transform 1 0 8800 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_340
timestamp 1675432918
transform 1 0 9350 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_341
timestamp 1675432918
transform 1 0 9350 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_342
timestamp 1675432918
transform 1 0 9350 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_343
timestamp 1675432918
transform 1 0 9350 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_344
timestamp 1675432918
transform 1 0 9350 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_345
timestamp 1675432918
transform 1 0 9350 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_346
timestamp 1675432918
transform 1 0 9350 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_347
timestamp 1675432918
transform 1 0 9350 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_348
timestamp 1675432918
transform 1 0 9350 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_349
timestamp 1675432918
transform 1 0 9350 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_350
timestamp 1675432918
transform 1 0 9350 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_351
timestamp 1675432918
transform 1 0 9350 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_352
timestamp 1675432918
transform 1 0 9350 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_353
timestamp 1675432918
transform 1 0 9350 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_354
timestamp 1675432918
transform 1 0 9350 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_355
timestamp 1675432918
transform 1 0 9350 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_356
timestamp 1675432918
transform 1 0 9350 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_357
timestamp 1675432918
transform 1 0 9350 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_358
timestamp 1675432918
transform 1 0 9350 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_359
timestamp 1675432918
transform 1 0 9350 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_360
timestamp 1675432918
transform 1 0 9900 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_361
timestamp 1675432918
transform 1 0 9900 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_362
timestamp 1675432918
transform 1 0 9900 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_363
timestamp 1675432918
transform 1 0 9900 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_364
timestamp 1675432918
transform 1 0 9900 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_365
timestamp 1675432918
transform 1 0 9900 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_366
timestamp 1675432918
transform 1 0 9900 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_367
timestamp 1675432918
transform 1 0 9900 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_368
timestamp 1675432918
transform 1 0 9900 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_369
timestamp 1675432918
transform 1 0 9900 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_370
timestamp 1675432918
transform 1 0 9900 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_371
timestamp 1675432918
transform 1 0 9900 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_372
timestamp 1675432918
transform 1 0 9900 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_373
timestamp 1675432918
transform 1 0 9900 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_374
timestamp 1675432918
transform 1 0 9900 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_375
timestamp 1675432918
transform 1 0 9900 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_376
timestamp 1675432918
transform 1 0 9900 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_377
timestamp 1675432918
transform 1 0 9900 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_378
timestamp 1675432918
transform 1 0 9900 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_379
timestamp 1675432918
transform 1 0 9900 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_380
timestamp 1675432918
transform 1 0 10450 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_381
timestamp 1675432918
transform 1 0 10450 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_382
timestamp 1675432918
transform 1 0 10450 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_383
timestamp 1675432918
transform 1 0 10450 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_384
timestamp 1675432918
transform 1 0 10450 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_385
timestamp 1675432918
transform 1 0 10450 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_386
timestamp 1675432918
transform 1 0 10450 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_387
timestamp 1675432918
transform 1 0 10450 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_388
timestamp 1675432918
transform 1 0 10450 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_389
timestamp 1675432918
transform 1 0 10450 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_390
timestamp 1675432918
transform 1 0 10450 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_391
timestamp 1675432918
transform 1 0 10450 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_392
timestamp 1675432918
transform 1 0 10450 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_393
timestamp 1675432918
transform 1 0 10450 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_394
timestamp 1675432918
transform 1 0 10450 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_395
timestamp 1675432918
transform 1 0 10450 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_396
timestamp 1675432918
transform 1 0 10450 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_397
timestamp 1675432918
transform 1 0 10450 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_398
timestamp 1675432918
transform 1 0 10450 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_399
timestamp 1675432918
transform 1 0 10450 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_400
timestamp 1675432918
transform 1 0 11000 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_401
timestamp 1675432918
transform 1 0 11000 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_402
timestamp 1675432918
transform 1 0 11000 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_403
timestamp 1675432918
transform 1 0 11000 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_404
timestamp 1675432918
transform 1 0 11000 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_405
timestamp 1675432918
transform 1 0 11000 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_406
timestamp 1675432918
transform 1 0 11000 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_407
timestamp 1675432918
transform 1 0 11000 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_408
timestamp 1675432918
transform 1 0 11000 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_409
timestamp 1675432918
transform 1 0 11000 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_410
timestamp 1675432918
transform 1 0 11000 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_411
timestamp 1675432918
transform 1 0 11000 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_412
timestamp 1675432918
transform 1 0 11000 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_413
timestamp 1675432918
transform 1 0 11000 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_414
timestamp 1675432918
transform 1 0 11000 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_415
timestamp 1675432918
transform 1 0 11000 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_416
timestamp 1675432918
transform 1 0 11000 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_417
timestamp 1675432918
transform 1 0 11000 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_418
timestamp 1675432918
transform 1 0 11000 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_419
timestamp 1675432918
transform 1 0 11000 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_420
timestamp 1675432918
transform 1 0 11550 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_421
timestamp 1675432918
transform 1 0 11550 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_422
timestamp 1675432918
transform 1 0 11550 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_423
timestamp 1675432918
transform 1 0 11550 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_424
timestamp 1675432918
transform 1 0 11550 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_425
timestamp 1675432918
transform 1 0 11550 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_426
timestamp 1675432918
transform 1 0 11550 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_427
timestamp 1675432918
transform 1 0 11550 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_428
timestamp 1675432918
transform 1 0 11550 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_429
timestamp 1675432918
transform 1 0 11550 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_430
timestamp 1675432918
transform 1 0 11550 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_431
timestamp 1675432918
transform 1 0 11550 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_432
timestamp 1675432918
transform 1 0 11550 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_433
timestamp 1675432918
transform 1 0 11550 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_434
timestamp 1675432918
transform 1 0 11550 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_435
timestamp 1675432918
transform 1 0 11550 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_436
timestamp 1675432918
transform 1 0 11550 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_437
timestamp 1675432918
transform 1 0 11550 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_438
timestamp 1675432918
transform 1 0 11550 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_439
timestamp 1675432918
transform 1 0 11550 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_440
timestamp 1675432918
transform 1 0 12100 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_441
timestamp 1675432918
transform 1 0 12100 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_442
timestamp 1675432918
transform 1 0 12100 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_443
timestamp 1675432918
transform 1 0 12100 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_444
timestamp 1675432918
transform 1 0 12100 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_445
timestamp 1675432918
transform 1 0 12100 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_446
timestamp 1675432918
transform 1 0 12100 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_447
timestamp 1675432918
transform 1 0 12100 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_448
timestamp 1675432918
transform 1 0 12100 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_449
timestamp 1675432918
transform 1 0 12100 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_450
timestamp 1675432918
transform 1 0 12100 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_451
timestamp 1675432918
transform 1 0 12100 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_452
timestamp 1675432918
transform 1 0 12100 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_453
timestamp 1675432918
transform 1 0 12100 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_454
timestamp 1675432918
transform 1 0 12100 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_455
timestamp 1675432918
transform 1 0 12100 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_456
timestamp 1675432918
transform 1 0 12100 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_457
timestamp 1675432918
transform 1 0 12100 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_458
timestamp 1675432918
transform 1 0 12100 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_459
timestamp 1675432918
transform 1 0 12100 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_460
timestamp 1675432918
transform 1 0 12650 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_461
timestamp 1675432918
transform 1 0 12650 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_462
timestamp 1675432918
transform 1 0 12650 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_463
timestamp 1675432918
transform 1 0 12650 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_464
timestamp 1675432918
transform 1 0 12650 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_465
timestamp 1675432918
transform 1 0 12650 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_466
timestamp 1675432918
transform 1 0 12650 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_467
timestamp 1675432918
transform 1 0 12650 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_468
timestamp 1675432918
transform 1 0 12650 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_469
timestamp 1675432918
transform 1 0 12650 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_470
timestamp 1675432918
transform 1 0 12650 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_471
timestamp 1675432918
transform 1 0 12650 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_472
timestamp 1675432918
transform 1 0 12650 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_473
timestamp 1675432918
transform 1 0 12650 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_474
timestamp 1675432918
transform 1 0 12650 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_475
timestamp 1675432918
transform 1 0 12650 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_476
timestamp 1675432918
transform 1 0 12650 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_477
timestamp 1675432918
transform 1 0 12650 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_478
timestamp 1675432918
transform 1 0 12650 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_479
timestamp 1675432918
transform 1 0 12650 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_480
timestamp 1675432918
transform 1 0 13200 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_481
timestamp 1675432918
transform 1 0 13200 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_482
timestamp 1675432918
transform 1 0 13200 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_483
timestamp 1675432918
transform 1 0 13200 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_484
timestamp 1675432918
transform 1 0 13200 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_485
timestamp 1675432918
transform 1 0 13200 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_486
timestamp 1675432918
transform 1 0 13200 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_487
timestamp 1675432918
transform 1 0 13200 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_488
timestamp 1675432918
transform 1 0 13200 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_489
timestamp 1675432918
transform 1 0 13200 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_490
timestamp 1675432918
transform 1 0 13200 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_491
timestamp 1675432918
transform 1 0 13200 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_492
timestamp 1675432918
transform 1 0 13200 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_493
timestamp 1675432918
transform 1 0 13200 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_494
timestamp 1675432918
transform 1 0 13200 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_495
timestamp 1675432918
transform 1 0 13200 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_496
timestamp 1675432918
transform 1 0 13200 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_497
timestamp 1675432918
transform 1 0 13200 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_498
timestamp 1675432918
transform 1 0 13200 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_499
timestamp 1675432918
transform 1 0 13200 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_500
timestamp 1675432918
transform 1 0 13750 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_501
timestamp 1675432918
transform 1 0 13750 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_502
timestamp 1675432918
transform 1 0 13750 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_503
timestamp 1675432918
transform 1 0 13750 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_504
timestamp 1675432918
transform 1 0 13750 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_505
timestamp 1675432918
transform 1 0 13750 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_506
timestamp 1675432918
transform 1 0 13750 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_507
timestamp 1675432918
transform 1 0 13750 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_508
timestamp 1675432918
transform 1 0 13750 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_509
timestamp 1675432918
transform 1 0 13750 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_510
timestamp 1675432918
transform 1 0 13750 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_511
timestamp 1675432918
transform 1 0 13750 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_512
timestamp 1675432918
transform 1 0 13750 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_513
timestamp 1675432918
transform 1 0 13750 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_514
timestamp 1675432918
transform 1 0 13750 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_515
timestamp 1675432918
transform 1 0 13750 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_516
timestamp 1675432918
transform 1 0 13750 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_517
timestamp 1675432918
transform 1 0 13750 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_518
timestamp 1675432918
transform 1 0 13750 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_519
timestamp 1675432918
transform 1 0 13750 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_520
timestamp 1675432918
transform 1 0 14300 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_521
timestamp 1675432918
transform 1 0 14300 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_522
timestamp 1675432918
transform 1 0 14300 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_523
timestamp 1675432918
transform 1 0 14300 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_524
timestamp 1675432918
transform 1 0 14300 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_525
timestamp 1675432918
transform 1 0 14300 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_526
timestamp 1675432918
transform 1 0 14300 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_527
timestamp 1675432918
transform 1 0 14300 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_528
timestamp 1675432918
transform 1 0 14300 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_529
timestamp 1675432918
transform 1 0 14300 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_530
timestamp 1675432918
transform 1 0 14300 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_531
timestamp 1675432918
transform 1 0 14300 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_532
timestamp 1675432918
transform 1 0 14300 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_533
timestamp 1675432918
transform 1 0 14300 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_534
timestamp 1675432918
transform 1 0 14300 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_535
timestamp 1675432918
transform 1 0 14300 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_536
timestamp 1675432918
transform 1 0 14300 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_537
timestamp 1675432918
transform 1 0 14300 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_538
timestamp 1675432918
transform 1 0 14300 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_539
timestamp 1675432918
transform 1 0 14300 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_540
timestamp 1675432918
transform 1 0 14850 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_541
timestamp 1675432918
transform 1 0 14850 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_542
timestamp 1675432918
transform 1 0 14850 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_543
timestamp 1675432918
transform 1 0 14850 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_544
timestamp 1675432918
transform 1 0 14850 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_545
timestamp 1675432918
transform 1 0 14850 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_546
timestamp 1675432918
transform 1 0 14850 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_547
timestamp 1675432918
transform 1 0 14850 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_548
timestamp 1675432918
transform 1 0 14850 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_549
timestamp 1675432918
transform 1 0 14850 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_550
timestamp 1675432918
transform 1 0 14850 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_551
timestamp 1675432918
transform 1 0 14850 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_552
timestamp 1675432918
transform 1 0 14850 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_553
timestamp 1675432918
transform 1 0 14850 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_554
timestamp 1675432918
transform 1 0 14850 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_555
timestamp 1675432918
transform 1 0 14850 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_556
timestamp 1675432918
transform 1 0 14850 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_557
timestamp 1675432918
transform 1 0 14850 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_558
timestamp 1675432918
transform 1 0 14850 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_559
timestamp 1675432918
transform 1 0 14850 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_560
timestamp 1675432918
transform 1 0 15400 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_561
timestamp 1675432918
transform 1 0 15400 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_562
timestamp 1675432918
transform 1 0 15400 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_563
timestamp 1675432918
transform 1 0 15400 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_564
timestamp 1675432918
transform 1 0 15400 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_565
timestamp 1675432918
transform 1 0 15400 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_566
timestamp 1675432918
transform 1 0 15400 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_567
timestamp 1675432918
transform 1 0 15400 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_568
timestamp 1675432918
transform 1 0 15400 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_569
timestamp 1675432918
transform 1 0 15400 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_570
timestamp 1675432918
transform 1 0 15400 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_571
timestamp 1675432918
transform 1 0 15400 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_572
timestamp 1675432918
transform 1 0 15400 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_573
timestamp 1675432918
transform 1 0 15400 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_574
timestamp 1675432918
transform 1 0 15400 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_575
timestamp 1675432918
transform 1 0 15400 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_576
timestamp 1675432918
transform 1 0 15400 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_577
timestamp 1675432918
transform 1 0 15400 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_578
timestamp 1675432918
transform 1 0 15400 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_579
timestamp 1675432918
transform 1 0 15400 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_580
timestamp 1675432918
transform 1 0 15950 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_581
timestamp 1675432918
transform 1 0 15950 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_582
timestamp 1675432918
transform 1 0 15950 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_583
timestamp 1675432918
transform 1 0 15950 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_584
timestamp 1675432918
transform 1 0 15950 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_585
timestamp 1675432918
transform 1 0 15950 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_586
timestamp 1675432918
transform 1 0 15950 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_587
timestamp 1675432918
transform 1 0 15950 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_588
timestamp 1675432918
transform 1 0 15950 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_589
timestamp 1675432918
transform 1 0 15950 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_590
timestamp 1675432918
transform 1 0 15950 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_591
timestamp 1675432918
transform 1 0 15950 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_592
timestamp 1675432918
transform 1 0 15950 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_593
timestamp 1675432918
transform 1 0 15950 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_594
timestamp 1675432918
transform 1 0 15950 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_595
timestamp 1675432918
transform 1 0 15950 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_596
timestamp 1675432918
transform 1 0 15950 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_597
timestamp 1675432918
transform 1 0 15950 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_598
timestamp 1675432918
transform 1 0 15950 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_599
timestamp 1675432918
transform 1 0 15950 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_600
timestamp 1675432918
transform 1 0 16500 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_601
timestamp 1675432918
transform 1 0 16500 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_602
timestamp 1675432918
transform 1 0 16500 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_603
timestamp 1675432918
transform 1 0 16500 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_604
timestamp 1675432918
transform 1 0 16500 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_605
timestamp 1675432918
transform 1 0 16500 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_606
timestamp 1675432918
transform 1 0 16500 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_607
timestamp 1675432918
transform 1 0 16500 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_608
timestamp 1675432918
transform 1 0 16500 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_609
timestamp 1675432918
transform 1 0 16500 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_610
timestamp 1675432918
transform 1 0 16500 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_611
timestamp 1675432918
transform 1 0 16500 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_612
timestamp 1675432918
transform 1 0 16500 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_613
timestamp 1675432918
transform 1 0 16500 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_614
timestamp 1675432918
transform 1 0 16500 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_615
timestamp 1675432918
transform 1 0 16500 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_616
timestamp 1675432918
transform 1 0 16500 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_617
timestamp 1675432918
transform 1 0 16500 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_618
timestamp 1675432918
transform 1 0 16500 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_619
timestamp 1675432918
transform 1 0 16500 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_620
timestamp 1675432918
transform 1 0 17050 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_621
timestamp 1675432918
transform 1 0 17050 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_622
timestamp 1675432918
transform 1 0 17050 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_623
timestamp 1675432918
transform 1 0 17050 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_624
timestamp 1675432918
transform 1 0 17050 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_625
timestamp 1675432918
transform 1 0 17050 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_626
timestamp 1675432918
transform 1 0 17050 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_627
timestamp 1675432918
transform 1 0 17050 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_628
timestamp 1675432918
transform 1 0 17050 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_629
timestamp 1675432918
transform 1 0 17050 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_630
timestamp 1675432918
transform 1 0 17050 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_631
timestamp 1675432918
transform 1 0 17050 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_632
timestamp 1675432918
transform 1 0 17050 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_633
timestamp 1675432918
transform 1 0 17050 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_634
timestamp 1675432918
transform 1 0 17050 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_635
timestamp 1675432918
transform 1 0 17050 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_636
timestamp 1675432918
transform 1 0 17050 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_637
timestamp 1675432918
transform 1 0 17050 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_638
timestamp 1675432918
transform 1 0 17050 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_639
timestamp 1675432918
transform 1 0 17050 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_640
timestamp 1675432918
transform 1 0 17600 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_641
timestamp 1675432918
transform 1 0 17600 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_642
timestamp 1675432918
transform 1 0 17600 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_643
timestamp 1675432918
transform 1 0 17600 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_644
timestamp 1675432918
transform 1 0 17600 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_645
timestamp 1675432918
transform 1 0 17600 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_646
timestamp 1675432918
transform 1 0 17600 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_647
timestamp 1675432918
transform 1 0 17600 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_648
timestamp 1675432918
transform 1 0 17600 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_649
timestamp 1675432918
transform 1 0 17600 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_650
timestamp 1675432918
transform 1 0 17600 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_651
timestamp 1675432918
transform 1 0 17600 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_652
timestamp 1675432918
transform 1 0 17600 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_653
timestamp 1675432918
transform 1 0 17600 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_654
timestamp 1675432918
transform 1 0 17600 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_655
timestamp 1675432918
transform 1 0 17600 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_656
timestamp 1675432918
transform 1 0 17600 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_657
timestamp 1675432918
transform 1 0 17600 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_658
timestamp 1675432918
transform 1 0 17600 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_659
timestamp 1675432918
transform 1 0 17600 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_660
timestamp 1675432918
transform 1 0 18150 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_661
timestamp 1675432918
transform 1 0 18150 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_662
timestamp 1675432918
transform 1 0 18150 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_663
timestamp 1675432918
transform 1 0 18150 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_664
timestamp 1675432918
transform 1 0 18150 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_665
timestamp 1675432918
transform 1 0 18150 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_666
timestamp 1675432918
transform 1 0 18150 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_667
timestamp 1675432918
transform 1 0 18150 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_668
timestamp 1675432918
transform 1 0 18150 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_669
timestamp 1675432918
transform 1 0 18150 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_670
timestamp 1675432918
transform 1 0 18150 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_671
timestamp 1675432918
transform 1 0 18150 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_672
timestamp 1675432918
transform 1 0 18150 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_673
timestamp 1675432918
transform 1 0 18150 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_674
timestamp 1675432918
transform 1 0 18150 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_675
timestamp 1675432918
transform 1 0 18150 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_676
timestamp 1675432918
transform 1 0 18150 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_677
timestamp 1675432918
transform 1 0 18150 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_678
timestamp 1675432918
transform 1 0 18150 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_679
timestamp 1675432918
transform 1 0 18150 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_680
timestamp 1675432918
transform 1 0 18700 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_681
timestamp 1675432918
transform 1 0 18700 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_682
timestamp 1675432918
transform 1 0 18700 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_683
timestamp 1675432918
transform 1 0 18700 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_684
timestamp 1675432918
transform 1 0 18700 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_685
timestamp 1675432918
transform 1 0 18700 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_686
timestamp 1675432918
transform 1 0 18700 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_687
timestamp 1675432918
transform 1 0 18700 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_688
timestamp 1675432918
transform 1 0 18700 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_689
timestamp 1675432918
transform 1 0 18700 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_690
timestamp 1675432918
transform 1 0 18700 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_691
timestamp 1675432918
transform 1 0 18700 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_692
timestamp 1675432918
transform 1 0 18700 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_693
timestamp 1675432918
transform 1 0 18700 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_694
timestamp 1675432918
transform 1 0 18700 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_695
timestamp 1675432918
transform 1 0 18700 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_696
timestamp 1675432918
transform 1 0 18700 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_697
timestamp 1675432918
transform 1 0 18700 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_698
timestamp 1675432918
transform 1 0 18700 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_699
timestamp 1675432918
transform 1 0 18700 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_700
timestamp 1675432918
transform 1 0 19250 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_701
timestamp 1675432918
transform 1 0 19250 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_702
timestamp 1675432918
transform 1 0 19250 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_703
timestamp 1675432918
transform 1 0 19250 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_704
timestamp 1675432918
transform 1 0 19250 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_705
timestamp 1675432918
transform 1 0 19250 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_706
timestamp 1675432918
transform 1 0 19250 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_707
timestamp 1675432918
transform 1 0 19250 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_708
timestamp 1675432918
transform 1 0 19250 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_709
timestamp 1675432918
transform 1 0 19250 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_710
timestamp 1675432918
transform 1 0 19250 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_711
timestamp 1675432918
transform 1 0 19250 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_712
timestamp 1675432918
transform 1 0 19250 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_713
timestamp 1675432918
transform 1 0 19250 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_714
timestamp 1675432918
transform 1 0 19250 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_715
timestamp 1675432918
transform 1 0 19250 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_716
timestamp 1675432918
transform 1 0 19250 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_717
timestamp 1675432918
transform 1 0 19250 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_718
timestamp 1675432918
transform 1 0 19250 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_719
timestamp 1675432918
transform 1 0 19250 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_720
timestamp 1675432918
transform 1 0 19800 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_721
timestamp 1675432918
transform 1 0 19800 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_722
timestamp 1675432918
transform 1 0 19800 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_723
timestamp 1675432918
transform 1 0 19800 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_724
timestamp 1675432918
transform 1 0 19800 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_725
timestamp 1675432918
transform 1 0 19800 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_726
timestamp 1675432918
transform 1 0 19800 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_727
timestamp 1675432918
transform 1 0 19800 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_728
timestamp 1675432918
transform 1 0 19800 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_729
timestamp 1675432918
transform 1 0 19800 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_730
timestamp 1675432918
transform 1 0 19800 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_731
timestamp 1675432918
transform 1 0 19800 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_732
timestamp 1675432918
transform 1 0 19800 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_733
timestamp 1675432918
transform 1 0 19800 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_734
timestamp 1675432918
transform 1 0 19800 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_735
timestamp 1675432918
transform 1 0 19800 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_736
timestamp 1675432918
transform 1 0 19800 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_737
timestamp 1675432918
transform 1 0 19800 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_738
timestamp 1675432918
transform 1 0 19800 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_739
timestamp 1675432918
transform 1 0 19800 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_740
timestamp 1675432918
transform 1 0 20350 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_741
timestamp 1675432918
transform 1 0 20350 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_742
timestamp 1675432918
transform 1 0 20350 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_743
timestamp 1675432918
transform 1 0 20350 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_744
timestamp 1675432918
transform 1 0 20350 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_745
timestamp 1675432918
transform 1 0 20350 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_746
timestamp 1675432918
transform 1 0 20350 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_747
timestamp 1675432918
transform 1 0 20350 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_748
timestamp 1675432918
transform 1 0 20350 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_749
timestamp 1675432918
transform 1 0 20350 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_750
timestamp 1675432918
transform 1 0 20350 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_751
timestamp 1675432918
transform 1 0 20350 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_752
timestamp 1675432918
transform 1 0 20350 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_753
timestamp 1675432918
transform 1 0 20350 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_754
timestamp 1675432918
transform 1 0 20350 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_755
timestamp 1675432918
transform 1 0 20350 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_756
timestamp 1675432918
transform 1 0 20350 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_757
timestamp 1675432918
transform 1 0 20350 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_758
timestamp 1675432918
transform 1 0 20350 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_759
timestamp 1675432918
transform 1 0 20350 0 1 21450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_760
timestamp 1675432918
transform 1 0 20900 0 1 0
box -113 -113 663 663
use pmos_source_in  pmos_source_in_761
timestamp 1675432918
transform 1 0 20900 0 1 1100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_762
timestamp 1675432918
transform 1 0 20900 0 1 2200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_763
timestamp 1675432918
transform 1 0 20900 0 1 3300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_764
timestamp 1675432918
transform 1 0 20900 0 1 4400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_765
timestamp 1675432918
transform 1 0 20900 0 1 5500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_766
timestamp 1675432918
transform 1 0 20900 0 1 6600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_767
timestamp 1675432918
transform 1 0 20900 0 1 7700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_768
timestamp 1675432918
transform 1 0 20900 0 1 8800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_769
timestamp 1675432918
transform 1 0 20900 0 1 9900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_770
timestamp 1675432918
transform 1 0 20900 0 1 11000
box -113 -113 663 663
use pmos_source_in  pmos_source_in_771
timestamp 1675432918
transform 1 0 20900 0 1 12100
box -113 -113 663 663
use pmos_source_in  pmos_source_in_772
timestamp 1675432918
transform 1 0 20900 0 1 13200
box -113 -113 663 663
use pmos_source_in  pmos_source_in_773
timestamp 1675432918
transform 1 0 20900 0 1 14300
box -113 -113 663 663
use pmos_source_in  pmos_source_in_774
timestamp 1675432918
transform 1 0 20900 0 1 15400
box -113 -113 663 663
use pmos_source_in  pmos_source_in_775
timestamp 1675432918
transform 1 0 20900 0 1 16500
box -113 -113 663 663
use pmos_source_in  pmos_source_in_776
timestamp 1675432918
transform 1 0 20900 0 1 17600
box -113 -113 663 663
use pmos_source_in  pmos_source_in_777
timestamp 1675432918
transform 1 0 20900 0 1 18700
box -113 -113 663 663
use pmos_source_in  pmos_source_in_778
timestamp 1675432918
transform 1 0 20900 0 1 19800
box -113 -113 663 663
use pmos_source_in  pmos_source_in_779
timestamp 1675432918
transform 1 0 20900 0 1 20900
box -113 -113 663 663
use pmos_source_in  pmos_source_in_780
timestamp 1675432918
transform 1 0 21450 0 1 550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_781
timestamp 1675432918
transform 1 0 21450 0 1 1650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_782
timestamp 1675432918
transform 1 0 21450 0 1 2750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_783
timestamp 1675432918
transform 1 0 21450 0 1 3850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_784
timestamp 1675432918
transform 1 0 21450 0 1 4950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_785
timestamp 1675432918
transform 1 0 21450 0 1 6050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_786
timestamp 1675432918
transform 1 0 21450 0 1 7150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_787
timestamp 1675432918
transform 1 0 21450 0 1 8250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_788
timestamp 1675432918
transform 1 0 21450 0 1 9350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_789
timestamp 1675432918
transform 1 0 21450 0 1 10450
box -113 -113 663 663
use pmos_source_in  pmos_source_in_790
timestamp 1675432918
transform 1 0 21450 0 1 11550
box -113 -113 663 663
use pmos_source_in  pmos_source_in_791
timestamp 1675432918
transform 1 0 21450 0 1 12650
box -113 -113 663 663
use pmos_source_in  pmos_source_in_792
timestamp 1675432918
transform 1 0 21450 0 1 13750
box -113 -113 663 663
use pmos_source_in  pmos_source_in_793
timestamp 1675432918
transform 1 0 21450 0 1 14850
box -113 -113 663 663
use pmos_source_in  pmos_source_in_794
timestamp 1675432918
transform 1 0 21450 0 1 15950
box -113 -113 663 663
use pmos_source_in  pmos_source_in_795
timestamp 1675432918
transform 1 0 21450 0 1 17050
box -113 -113 663 663
use pmos_source_in  pmos_source_in_796
timestamp 1675432918
transform 1 0 21450 0 1 18150
box -113 -113 663 663
use pmos_source_in  pmos_source_in_797
timestamp 1675432918
transform 1 0 21450 0 1 19250
box -113 -113 663 663
use pmos_source_in  pmos_source_in_798
timestamp 1675432918
transform 1 0 21450 0 1 20350
box -113 -113 663 663
use pmos_source_in  pmos_source_in_799
timestamp 1675432918
transform 1 0 21450 0 1 21450
box -113 -113 663 663
<< end >>
