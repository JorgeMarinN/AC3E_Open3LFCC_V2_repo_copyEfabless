magic
tech sky130A
magscale 1 2
timestamp 1699804740
<< checkpaint >>
rect -2866 -1804 30834 31724
<< viali >>
rect 3893 27557 3927 27591
rect 10609 27557 10643 27591
rect 17785 27557 17819 27591
rect 24869 27557 24903 27591
rect 4169 27353 4203 27387
rect 6929 27353 6963 27387
rect 7113 27353 7147 27387
rect 10885 27353 10919 27387
rect 17601 27353 17635 27387
rect 24593 27353 24627 27387
rect 6745 27285 6779 27319
rect 4261 27081 4295 27115
rect 6745 27013 6779 27047
rect 7573 27013 7607 27047
rect 4169 26945 4203 26979
rect 4445 26945 4479 26979
rect 4537 26945 4571 26979
rect 6561 26945 6595 26979
rect 6837 26945 6871 26979
rect 6929 26945 6963 26979
rect 7205 26945 7239 26979
rect 7389 26945 7423 26979
rect 10241 26945 10275 26979
rect 10977 26945 11011 26979
rect 12633 26945 12667 26979
rect 13185 26945 13219 26979
rect 17325 26945 17359 26979
rect 17417 26945 17451 26979
rect 5181 26877 5215 26911
rect 19717 26877 19751 26911
rect 19993 26877 20027 26911
rect 4445 26741 4479 26775
rect 7113 26741 7147 26775
rect 10333 26741 10367 26775
rect 11069 26741 11103 26775
rect 12725 26741 12759 26775
rect 13093 26741 13127 26775
rect 16681 26741 16715 26775
rect 17509 26741 17543 26775
rect 18245 26741 18279 26775
rect 6837 26537 6871 26571
rect 14427 26537 14461 26571
rect 15991 26537 16025 26571
rect 18981 26537 19015 26571
rect 3617 26469 3651 26503
rect 8677 26469 8711 26503
rect 15853 26469 15887 26503
rect 4077 26401 4111 26435
rect 6561 26401 6595 26435
rect 6929 26401 6963 26435
rect 17785 26401 17819 26435
rect 19257 26401 19291 26435
rect 26157 26401 26191 26435
rect 3341 26333 3375 26367
rect 3617 26333 3651 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4445 26333 4479 26367
rect 6469 26333 6503 26367
rect 7297 26333 7331 26367
rect 9045 26333 9079 26367
rect 9137 26333 9171 26367
rect 10885 26333 10919 26367
rect 11253 26333 11287 26367
rect 11345 26333 11379 26367
rect 13553 26333 13587 26367
rect 13737 26333 13771 26367
rect 13921 26333 13955 26367
rect 14105 26333 14139 26367
rect 14289 26333 14323 26367
rect 14565 26333 14599 26367
rect 14841 26333 14875 26367
rect 15577 26333 15611 26367
rect 17417 26333 17451 26367
rect 18061 26333 18095 26367
rect 18889 26333 18923 26367
rect 25513 26333 25547 26367
rect 5871 26265 5905 26299
rect 9413 26265 9447 26299
rect 11621 26265 11655 26299
rect 13645 26265 13679 26299
rect 15853 26265 15887 26299
rect 19533 26265 19567 26299
rect 21281 26265 21315 26299
rect 3433 26197 3467 26231
rect 3893 26197 3927 26231
rect 13093 26197 13127 26231
rect 13369 26197 13403 26231
rect 14105 26197 14139 26231
rect 14749 26197 14783 26231
rect 15669 26197 15703 26231
rect 17969 26197 18003 26231
rect 5089 25993 5123 26027
rect 7297 25993 7331 26027
rect 11345 25993 11379 26027
rect 18475 25993 18509 26027
rect 19625 25993 19659 26027
rect 4813 25925 4847 25959
rect 11989 25925 12023 25959
rect 12127 25925 12161 25959
rect 16313 25925 16347 25959
rect 2789 25857 2823 25891
rect 3157 25857 3191 25891
rect 4905 25857 4939 25891
rect 4997 25857 5031 25891
rect 7021 25857 7055 25891
rect 7481 25857 7515 25891
rect 7757 25857 7791 25891
rect 7941 25857 7975 25891
rect 10425 25857 10459 25891
rect 11069 25857 11103 25891
rect 11805 25857 11839 25891
rect 11897 25857 11931 25891
rect 12265 25857 12299 25891
rect 12357 25857 12391 25891
rect 12541 25857 12575 25891
rect 15761 25857 15795 25891
rect 15945 25857 15979 25891
rect 16037 25857 16071 25891
rect 16129 25857 16163 25891
rect 17049 25857 17083 25891
rect 19533 25857 19567 25891
rect 7113 25789 7147 25823
rect 7665 25789 7699 25823
rect 8631 25789 8665 25823
rect 10057 25789 10091 25823
rect 10885 25789 10919 25823
rect 10977 25789 11011 25823
rect 11161 25789 11195 25823
rect 12633 25789 12667 25823
rect 13369 25789 13403 25823
rect 13737 25789 13771 25823
rect 16681 25789 16715 25823
rect 7757 25721 7791 25755
rect 12449 25721 12483 25755
rect 15945 25721 15979 25755
rect 4583 25653 4617 25687
rect 6653 25653 6687 25687
rect 11621 25653 11655 25687
rect 13277 25653 13311 25687
rect 15163 25653 15197 25687
rect 16313 25653 16347 25687
rect 4629 25449 4663 25483
rect 7113 25449 7147 25483
rect 9965 25449 9999 25483
rect 11529 25449 11563 25483
rect 12265 25449 12299 25483
rect 13921 25449 13955 25483
rect 15485 25449 15519 25483
rect 19809 25449 19843 25483
rect 4445 25381 4479 25415
rect 11437 25381 11471 25415
rect 12633 25381 12667 25415
rect 13461 25381 13495 25415
rect 4077 25313 4111 25347
rect 9781 25313 9815 25347
rect 11161 25313 11195 25347
rect 11897 25313 11931 25347
rect 13829 25313 13863 25347
rect 14381 25313 14415 25347
rect 14933 25313 14967 25347
rect 15669 25313 15703 25347
rect 16129 25313 16163 25347
rect 18613 25313 18647 25347
rect 3985 25245 4019 25279
rect 4905 25245 4939 25279
rect 6837 25245 6871 25279
rect 9137 25245 9171 25279
rect 10057 25245 10091 25279
rect 10149 25245 10183 25279
rect 11069 25245 11103 25279
rect 11713 25245 11747 25279
rect 11805 25245 11839 25279
rect 11989 25245 12023 25279
rect 12449 25245 12483 25279
rect 12541 25245 12575 25279
rect 12725 25245 12759 25279
rect 13645 25245 13679 25279
rect 14289 25245 14323 25279
rect 14473 25245 14507 25279
rect 14565 25245 14599 25279
rect 14841 25245 14875 25279
rect 15025 25245 15059 25279
rect 15301 25245 15335 25279
rect 15761 25245 15795 25279
rect 16221 25245 16255 25279
rect 16589 25245 16623 25279
rect 18521 25245 18555 25279
rect 19349 25245 19383 25279
rect 19441 25245 19475 25279
rect 19533 25245 19567 25279
rect 19625 25245 19659 25279
rect 4813 25177 4847 25211
rect 7097 25177 7131 25211
rect 7297 25177 7331 25211
rect 13921 25177 13955 25211
rect 15117 25177 15151 25211
rect 16405 25177 16439 25211
rect 16497 25177 16531 25211
rect 4353 25109 4387 25143
rect 4613 25109 4647 25143
rect 4997 25109 5031 25143
rect 6745 25109 6779 25143
rect 6929 25109 6963 25143
rect 10241 25109 10275 25143
rect 14105 25109 14139 25143
rect 16773 25109 16807 25143
rect 18889 25109 18923 25143
rect 4537 24905 4571 24939
rect 11897 24905 11931 24939
rect 12357 24905 12391 24939
rect 16129 24905 16163 24939
rect 4261 24837 4295 24871
rect 12081 24837 12115 24871
rect 13721 24837 13755 24871
rect 13921 24837 13955 24871
rect 15945 24837 15979 24871
rect 20177 24837 20211 24871
rect 1777 24769 1811 24803
rect 3985 24769 4019 24803
rect 4721 24769 4755 24803
rect 4813 24769 4847 24803
rect 4997 24769 5031 24803
rect 5457 24769 5491 24803
rect 6009 24769 6043 24803
rect 6193 24769 6227 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 6745 24769 6779 24803
rect 7389 24769 7423 24803
rect 7481 24769 7515 24803
rect 7665 24769 7699 24803
rect 7941 24769 7975 24803
rect 12265 24769 12299 24803
rect 12633 24769 12667 24803
rect 12909 24769 12943 24803
rect 13001 24769 13035 24803
rect 13093 24769 13127 24803
rect 13277 24769 13311 24803
rect 13461 24769 13495 24803
rect 15209 24769 15243 24803
rect 15761 24769 15795 24803
rect 18245 24769 18279 24803
rect 18521 24769 18555 24803
rect 18797 24769 18831 24803
rect 18955 24769 18989 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 19257 24769 19291 24803
rect 19441 24769 19475 24803
rect 20085 24769 20119 24803
rect 20361 24769 20395 24803
rect 2145 24701 2179 24735
rect 3893 24701 3927 24735
rect 4353 24701 4387 24735
rect 5365 24701 5399 24735
rect 5549 24701 5583 24735
rect 5641 24701 5675 24735
rect 6101 24701 6135 24735
rect 8033 24701 8067 24735
rect 8125 24701 8159 24735
rect 8217 24701 8251 24735
rect 15301 24701 15335 24735
rect 15577 24701 15611 24735
rect 18429 24701 18463 24735
rect 19809 24701 19843 24735
rect 20545 24701 20579 24735
rect 21833 24701 21867 24735
rect 22201 24701 22235 24735
rect 4905 24633 4939 24667
rect 7205 24633 7239 24667
rect 13553 24633 13587 24667
rect 18337 24633 18371 24667
rect 18705 24633 18739 24667
rect 19533 24633 19567 24667
rect 3571 24565 3605 24599
rect 3709 24565 3743 24599
rect 5181 24565 5215 24599
rect 6929 24565 6963 24599
rect 7665 24565 7699 24599
rect 7757 24565 7791 24599
rect 12541 24565 12575 24599
rect 13737 24565 13771 24599
rect 19717 24565 19751 24599
rect 23581 24565 23615 24599
rect 3433 24361 3467 24395
rect 4537 24361 4571 24395
rect 4721 24361 4755 24395
rect 6285 24361 6319 24395
rect 6975 24361 7009 24395
rect 7113 24361 7147 24395
rect 13185 24361 13219 24395
rect 13369 24361 13403 24395
rect 19257 24361 19291 24395
rect 22293 24361 22327 24395
rect 4077 24293 4111 24327
rect 7205 24293 7239 24327
rect 10333 24293 10367 24327
rect 19533 24293 19567 24327
rect 21557 24293 21591 24327
rect 1409 24225 1443 24259
rect 1777 24225 1811 24259
rect 19625 24225 19659 24259
rect 23305 24225 23339 24259
rect 3525 24157 3559 24191
rect 3985 24157 4019 24191
rect 4169 24157 4203 24191
rect 4261 24157 4295 24191
rect 4997 24157 5031 24191
rect 6469 24157 6503 24191
rect 6745 24157 6779 24191
rect 6837 24157 6871 24191
rect 7297 24157 7331 24191
rect 10057 24157 10091 24191
rect 13645 24157 13679 24191
rect 19441 24157 19475 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20085 24157 20119 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 22201 24157 22235 24191
rect 4675 24123 4709 24157
rect 3249 24089 3283 24123
rect 4905 24089 4939 24123
rect 5089 24089 5123 24123
rect 10333 24089 10367 24123
rect 13001 24089 13035 24123
rect 13201 24089 13235 24123
rect 4445 24021 4479 24055
rect 6653 24021 6687 24055
rect 10149 24021 10183 24055
rect 13553 24021 13587 24055
rect 22661 24021 22695 24055
rect 1593 23817 1627 23851
rect 2789 23817 2823 23851
rect 4169 23817 4203 23851
rect 8171 23817 8205 23851
rect 13553 23817 13587 23851
rect 19809 23817 19843 23851
rect 22477 23817 22511 23851
rect 2237 23749 2271 23783
rect 14657 23749 14691 23783
rect 19257 23749 19291 23783
rect 21649 23749 21683 23783
rect 19487 23715 19521 23749
rect 1409 23681 1443 23715
rect 2881 23681 2915 23715
rect 3893 23681 3927 23715
rect 3985 23681 4019 23715
rect 6377 23681 6411 23715
rect 6745 23681 6779 23715
rect 9229 23681 9263 23715
rect 9413 23681 9447 23715
rect 10308 23681 10342 23715
rect 10425 23681 10459 23715
rect 11345 23681 11379 23715
rect 13461 23681 13495 23715
rect 13645 23681 13679 23715
rect 13921 23681 13955 23715
rect 14381 23681 14415 23715
rect 16405 23681 16439 23715
rect 19717 23681 19751 23715
rect 21373 23681 21407 23715
rect 21465 23681 21499 23715
rect 21833 23681 21867 23715
rect 22017 23681 22051 23715
rect 22293 23681 22327 23715
rect 22569 23681 22603 23715
rect 22661 23681 22695 23715
rect 4169 23613 4203 23647
rect 10149 23613 10183 23647
rect 11161 23613 11195 23647
rect 15209 23613 15243 23647
rect 9413 23545 9447 23579
rect 10701 23545 10735 23579
rect 19625 23545 19659 23579
rect 21649 23545 21683 23579
rect 2513 23477 2547 23511
rect 9505 23477 9539 23511
rect 13829 23477 13863 23511
rect 14473 23477 14507 23511
rect 16313 23477 16347 23511
rect 19441 23477 19475 23511
rect 22201 23477 22235 23511
rect 22293 23477 22327 23511
rect 22753 23477 22787 23511
rect 7113 23273 7147 23307
rect 8585 23273 8619 23307
rect 11713 23273 11747 23307
rect 12909 23273 12943 23307
rect 15485 23273 15519 23307
rect 18429 23273 18463 23307
rect 19901 23273 19935 23307
rect 20085 23273 20119 23307
rect 20913 23273 20947 23307
rect 12357 23205 12391 23239
rect 13369 23205 13403 23239
rect 3065 23137 3099 23171
rect 9597 23137 9631 23171
rect 9873 23137 9907 23171
rect 10149 23137 10183 23171
rect 10609 23137 10643 23171
rect 10793 23137 10827 23171
rect 11345 23137 11379 23171
rect 13277 23137 13311 23171
rect 17233 23137 17267 23171
rect 21925 23137 21959 23171
rect 2789 23069 2823 23103
rect 6285 23069 6319 23103
rect 7021 23069 7055 23103
rect 8217 23069 8251 23103
rect 9756 23069 9790 23103
rect 11069 23069 11103 23103
rect 11161 23069 11195 23103
rect 11437 23069 11471 23103
rect 12081 23069 12115 23103
rect 12357 23069 12391 23103
rect 12633 23069 12667 23103
rect 13645 23069 13679 23103
rect 16865 23069 16899 23103
rect 18337 23069 18371 23103
rect 18521 23069 18555 23103
rect 18797 23069 18831 23103
rect 19073 23069 19107 23103
rect 19257 23069 19291 23103
rect 19533 23069 19567 23103
rect 19671 23069 19705 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21373 23069 21407 23103
rect 21649 23069 21683 23103
rect 6009 23001 6043 23035
rect 8585 23001 8619 23035
rect 10885 23001 10919 23035
rect 12541 23001 12575 23035
rect 13369 23001 13403 23035
rect 18613 23001 18647 23035
rect 19441 23001 19475 23035
rect 20269 23001 20303 23035
rect 20563 23001 20597 23035
rect 20729 23001 20763 23035
rect 21281 23001 21315 23035
rect 8769 22933 8803 22967
rect 8953 22933 8987 22967
rect 11529 22933 11563 22967
rect 11713 22933 11747 22967
rect 12725 22933 12759 22967
rect 12909 22933 12943 22967
rect 13553 22933 13587 22967
rect 18981 22933 19015 22967
rect 19809 22933 19843 22967
rect 20069 22933 20103 22967
rect 21557 22933 21591 22967
rect 23397 22933 23431 22967
rect 9597 22729 9631 22763
rect 12817 22729 12851 22763
rect 15255 22729 15289 22763
rect 8769 22661 8803 22695
rect 22109 22661 22143 22695
rect 8401 22593 8435 22627
rect 9137 22593 9171 22627
rect 9413 22593 9447 22627
rect 9689 22593 9723 22627
rect 9965 22593 9999 22627
rect 10793 22593 10827 22627
rect 10977 22593 11011 22627
rect 11253 22593 11287 22627
rect 11713 22593 11747 22627
rect 11805 22593 11839 22627
rect 12081 22593 12115 22627
rect 12357 22593 12391 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 13093 22593 13127 22627
rect 13461 22593 13495 22627
rect 13829 22593 13863 22627
rect 15853 22593 15887 22627
rect 16681 22593 16715 22627
rect 20545 22593 20579 22627
rect 20637 22593 20671 22627
rect 20821 22593 20855 22627
rect 21097 22593 21131 22627
rect 21833 22593 21867 22627
rect 9229 22525 9263 22559
rect 9321 22525 9355 22559
rect 9781 22525 9815 22559
rect 11069 22525 11103 22559
rect 16129 22525 16163 22559
rect 16957 22525 16991 22559
rect 18705 22525 18739 22559
rect 18797 22525 18831 22559
rect 20269 22525 20303 22559
rect 21005 22525 21039 22559
rect 21465 22525 21499 22559
rect 23857 22525 23891 22559
rect 8953 22457 8987 22491
rect 10885 22457 10919 22491
rect 8769 22389 8803 22423
rect 9689 22389 9723 22423
rect 10149 22389 10183 22423
rect 10609 22389 10643 22423
rect 11529 22389 11563 22423
rect 11989 22389 12023 22423
rect 12173 22389 12207 22423
rect 13277 22389 13311 22423
rect 20637 22389 20671 22423
rect 4629 22185 4663 22219
rect 9137 22185 9171 22219
rect 9597 22185 9631 22219
rect 9965 22185 9999 22219
rect 11253 22185 11287 22219
rect 14197 22185 14231 22219
rect 18521 22185 18555 22219
rect 18981 22185 19015 22219
rect 19257 22185 19291 22219
rect 20545 22185 20579 22219
rect 21281 22185 21315 22219
rect 11529 22049 11563 22083
rect 11713 22049 11747 22083
rect 16497 22049 16531 22083
rect 17233 22049 17267 22083
rect 19533 22049 19567 22083
rect 19625 22049 19659 22083
rect 19718 22049 19752 22083
rect 20913 22049 20947 22083
rect 21557 22049 21591 22083
rect 22661 22049 22695 22083
rect 1409 21981 1443 22015
rect 2421 21981 2455 22015
rect 2881 21981 2915 22015
rect 3157 21981 3191 22015
rect 3249 21981 3283 22015
rect 3341 21981 3375 22015
rect 3433 21981 3467 22015
rect 3801 21981 3835 22015
rect 3985 21981 4019 22015
rect 4077 21981 4111 22015
rect 4169 21981 4203 22015
rect 4261 21981 4295 22015
rect 4905 21981 4939 22015
rect 5181 21981 5215 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 5917 21981 5951 22015
rect 9413 21981 9447 22015
rect 9597 21981 9631 22015
rect 11437 21981 11471 22015
rect 11621 21981 11655 22015
rect 12265 21981 12299 22015
rect 15945 21981 15979 22015
rect 16589 21981 16623 22015
rect 17141 21981 17175 22015
rect 18153 21981 18187 22015
rect 18705 21981 18739 22015
rect 18797 21981 18831 22015
rect 19441 21981 19475 22015
rect 20085 21981 20119 22015
rect 20729 21981 20763 22015
rect 21649 21981 21683 22015
rect 22569 21981 22603 22015
rect 4583 21947 4617 21981
rect 4813 21913 4847 21947
rect 6193 21913 6227 21947
rect 8953 21913 8987 21947
rect 9781 21913 9815 21947
rect 12081 21913 12115 21947
rect 15669 21913 15703 21947
rect 17509 21913 17543 21947
rect 18981 21913 19015 21947
rect 1593 21845 1627 21879
rect 2513 21845 2547 21879
rect 2789 21845 2823 21879
rect 2973 21845 3007 21879
rect 4445 21845 4479 21879
rect 4997 21845 5031 21879
rect 5273 21845 5307 21879
rect 5641 21845 5675 21879
rect 7665 21845 7699 21879
rect 9153 21845 9187 21879
rect 9321 21845 9355 21879
rect 9981 21845 10015 21879
rect 10149 21845 10183 21879
rect 11897 21845 11931 21879
rect 19993 21845 20027 21879
rect 4261 21641 4295 21675
rect 5549 21641 5583 21675
rect 6469 21641 6503 21675
rect 7113 21641 7147 21675
rect 14657 21641 14691 21675
rect 15301 21641 15335 21675
rect 15669 21641 15703 21675
rect 18245 21641 18279 21675
rect 3433 21573 3467 21607
rect 3893 21573 3927 21607
rect 6929 21573 6963 21607
rect 12265 21573 12299 21607
rect 1409 21505 1443 21539
rect 3683 21505 3717 21539
rect 3801 21505 3835 21539
rect 3985 21505 4019 21539
rect 4537 21505 4571 21539
rect 4813 21505 4847 21539
rect 4997 21505 5031 21539
rect 5181 21505 5215 21539
rect 5273 21505 5307 21539
rect 5365 21505 5399 21539
rect 6101 21505 6135 21539
rect 6653 21505 6687 21539
rect 7205 21505 7239 21539
rect 14289 21505 14323 21539
rect 14749 21505 14783 21539
rect 15393 21505 15427 21539
rect 15485 21505 15519 21539
rect 17785 21505 17819 21539
rect 18061 21505 18095 21539
rect 18245 21505 18279 21539
rect 1685 21437 1719 21471
rect 3525 21437 3559 21471
rect 5825 21437 5859 21471
rect 5917 21437 5951 21471
rect 6009 21437 6043 21471
rect 6745 21437 6779 21471
rect 14013 21437 14047 21471
rect 14565 21437 14599 21471
rect 4169 21369 4203 21403
rect 15117 21369 15151 21403
rect 4721 21301 4755 21335
rect 5641 21301 5675 21335
rect 6837 21301 6871 21335
rect 17923 21301 17957 21335
rect 3893 21097 3927 21131
rect 5181 21097 5215 21131
rect 13093 21097 13127 21131
rect 16957 21097 16991 21131
rect 3387 21029 3421 21063
rect 4261 21029 4295 21063
rect 13829 21029 13863 21063
rect 1593 20961 1627 20995
rect 1961 20961 1995 20995
rect 8953 20961 8987 20995
rect 9137 20961 9171 20995
rect 14565 20961 14599 20995
rect 14749 20961 14783 20995
rect 4077 20893 4111 20927
rect 4169 20893 4203 20927
rect 4353 20893 4387 20927
rect 4721 20893 4755 20927
rect 4813 20893 4847 20927
rect 4997 20893 5031 20927
rect 9229 20893 9263 20927
rect 10149 20893 10183 20927
rect 10241 20893 10275 20927
rect 10425 20893 10459 20927
rect 12909 20893 12943 20927
rect 13921 20893 13955 20927
rect 17509 20893 17543 20927
rect 7021 20825 7055 20859
rect 9965 20825 9999 20859
rect 14473 20825 14507 20859
rect 15669 20825 15703 20859
rect 5733 20757 5767 20791
rect 8953 20757 8987 20791
rect 9781 20757 9815 20791
rect 10241 20757 10275 20791
rect 14105 20757 14139 20791
rect 17601 20757 17635 20791
rect 3433 20553 3467 20587
rect 4077 20553 4111 20587
rect 4905 20553 4939 20587
rect 5549 20553 5583 20587
rect 8217 20553 8251 20587
rect 9137 20553 9171 20587
rect 9321 20553 9355 20587
rect 10885 20553 10919 20587
rect 3893 20485 3927 20519
rect 5165 20485 5199 20519
rect 5365 20485 5399 20519
rect 10149 20485 10183 20519
rect 11529 20485 11563 20519
rect 3065 20417 3099 20451
rect 3709 20417 3743 20451
rect 5457 20417 5491 20451
rect 5917 20417 5951 20451
rect 6469 20417 6503 20451
rect 8953 20417 8987 20451
rect 9939 20417 9973 20451
rect 10057 20417 10091 20451
rect 10241 20417 10275 20451
rect 10701 20417 10735 20451
rect 10977 20417 11011 20451
rect 11713 20417 11747 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 15945 20417 15979 20451
rect 16957 20417 16991 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 17325 20417 17359 20451
rect 19901 20417 19935 20451
rect 3157 20349 3191 20383
rect 4261 20349 4295 20383
rect 5641 20349 5675 20383
rect 6745 20349 6779 20383
rect 9781 20349 9815 20383
rect 15393 20349 15427 20383
rect 17417 20349 17451 20383
rect 18889 20349 18923 20383
rect 19165 20349 19199 20383
rect 4997 20281 5031 20315
rect 9689 20281 9723 20315
rect 10425 20281 10459 20315
rect 16405 20281 16439 20315
rect 5181 20213 5215 20247
rect 5779 20213 5813 20247
rect 8401 20213 8435 20247
rect 9321 20213 9355 20247
rect 10517 20213 10551 20247
rect 11897 20213 11931 20247
rect 16681 20213 16715 20247
rect 19993 20213 20027 20247
rect 6929 20009 6963 20043
rect 7297 20009 7331 20043
rect 9413 20009 9447 20043
rect 10977 20009 11011 20043
rect 11805 20009 11839 20043
rect 12173 20009 12207 20043
rect 16129 20009 16163 20043
rect 16497 20009 16531 20043
rect 18429 20009 18463 20043
rect 18705 20009 18739 20043
rect 14841 19941 14875 19975
rect 16037 19941 16071 19975
rect 17877 19941 17911 19975
rect 10793 19873 10827 19907
rect 14473 19873 14507 19907
rect 17325 19873 17359 19907
rect 1409 19805 1443 19839
rect 4997 19805 5031 19839
rect 5181 19805 5215 19839
rect 5365 19805 5399 19839
rect 5549 19805 5583 19839
rect 7021 19805 7055 19839
rect 7205 19805 7239 19839
rect 8493 19805 8527 19839
rect 8677 19805 8711 19839
rect 8769 19805 8803 19839
rect 9045 19805 9079 19839
rect 9781 19805 9815 19839
rect 10057 19805 10091 19839
rect 10333 19805 10367 19839
rect 10609 19805 10643 19839
rect 11069 19805 11103 19839
rect 11345 19805 11379 19839
rect 11437 19805 11471 19839
rect 11713 19805 11747 19839
rect 12265 19805 12299 19839
rect 12541 19805 12575 19839
rect 12725 19805 12759 19839
rect 14657 19805 14691 19839
rect 15393 19805 15427 19839
rect 15577 19805 15611 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 16221 19805 16255 19839
rect 16865 19805 16899 19839
rect 17049 19805 17083 19839
rect 17417 19805 17451 19839
rect 18153 19805 18187 19839
rect 18245 19805 18279 19839
rect 18797 19805 18831 19839
rect 18889 19805 18923 19839
rect 19257 19805 19291 19839
rect 4813 19737 4847 19771
rect 9413 19737 9447 19771
rect 9873 19737 9907 19771
rect 10793 19737 10827 19771
rect 11529 19737 11563 19771
rect 14933 19737 14967 19771
rect 15485 19737 15519 19771
rect 17509 19737 17543 19771
rect 19533 19737 19567 19771
rect 1593 19669 1627 19703
rect 4629 19669 4663 19703
rect 8309 19669 8343 19703
rect 9597 19669 9631 19703
rect 11161 19669 11195 19703
rect 12909 19669 12943 19703
rect 16957 19669 16991 19703
rect 17969 19669 18003 19703
rect 19073 19669 19107 19703
rect 21005 19669 21039 19703
rect 3347 19465 3381 19499
rect 3433 19465 3467 19499
rect 10333 19465 10367 19499
rect 11161 19465 11195 19499
rect 11713 19465 11747 19499
rect 14749 19465 14783 19499
rect 17049 19465 17083 19499
rect 20913 19465 20947 19499
rect 2513 19397 2547 19431
rect 5273 19397 5307 19431
rect 13737 19397 13771 19431
rect 15761 19397 15795 19431
rect 16681 19397 16715 19431
rect 2421 19329 2455 19363
rect 2789 19329 2823 19363
rect 2973 19329 3007 19363
rect 3065 19329 3099 19363
rect 3249 19329 3283 19363
rect 3525 19329 3559 19363
rect 3617 19329 3651 19363
rect 3801 19329 3835 19363
rect 4629 19329 4663 19363
rect 5089 19329 5123 19363
rect 5365 19329 5399 19363
rect 5457 19329 5491 19363
rect 5733 19329 5767 19363
rect 5917 19329 5951 19363
rect 6377 19329 6411 19363
rect 8769 19329 8803 19363
rect 9413 19329 9447 19363
rect 9505 19329 9539 19363
rect 9965 19329 9999 19363
rect 10517 19329 10551 19363
rect 10977 19329 11011 19363
rect 11069 19329 11103 19363
rect 11253 19329 11287 19363
rect 12173 19329 12207 19363
rect 14565 19329 14599 19363
rect 16129 19329 16163 19363
rect 16221 19329 16255 19363
rect 16497 19329 16531 19363
rect 16865 19329 16899 19363
rect 17325 19329 17359 19363
rect 19165 19329 19199 19363
rect 3709 19261 3743 19295
rect 4721 19261 4755 19295
rect 4997 19261 5031 19295
rect 6653 19261 6687 19295
rect 8401 19261 8435 19295
rect 9689 19261 9723 19295
rect 10701 19261 10735 19295
rect 10793 19261 10827 19295
rect 17601 19261 17635 19295
rect 19441 19261 19475 19295
rect 5641 19193 5675 19227
rect 10609 19193 10643 19227
rect 13921 19193 13955 19227
rect 15577 19193 15611 19227
rect 2789 19125 2823 19159
rect 6101 19125 6135 19159
rect 12081 19125 12115 19159
rect 19073 19125 19107 19159
rect 5089 18921 5123 18955
rect 6929 18921 6963 18955
rect 9597 18921 9631 18955
rect 9965 18921 9999 18955
rect 10977 18921 11011 18955
rect 12541 18921 12575 18955
rect 15577 18921 15611 18955
rect 17969 18921 18003 18955
rect 18889 18921 18923 18955
rect 20085 18921 20119 18955
rect 20453 18921 20487 18955
rect 10701 18853 10735 18887
rect 16681 18853 16715 18887
rect 19993 18853 20027 18887
rect 1777 18785 1811 18819
rect 3525 18785 3559 18819
rect 4629 18785 4663 18819
rect 5273 18785 5307 18819
rect 12909 18785 12943 18819
rect 14105 18785 14139 18819
rect 14381 18785 14415 18819
rect 17417 18785 17451 18819
rect 18521 18785 18555 18819
rect 19441 18785 19475 18819
rect 1501 18717 1535 18751
rect 3985 18717 4019 18751
rect 4721 18717 4755 18751
rect 5181 18717 5215 18751
rect 5365 18717 5399 18751
rect 6837 18717 6871 18751
rect 9137 18717 9171 18751
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 10517 18717 10551 18751
rect 10793 18717 10827 18751
rect 12449 18717 12483 18751
rect 15025 18717 15059 18751
rect 15117 18717 15151 18751
rect 15301 18717 15335 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 16037 18717 16071 18751
rect 16405 18717 16439 18751
rect 16589 18717 16623 18751
rect 17141 18717 17175 18751
rect 17601 18717 17635 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 18981 18717 19015 18751
rect 19533 18717 19567 18751
rect 20269 18717 20303 18751
rect 20361 18717 20395 18751
rect 26525 18717 26559 18751
rect 15853 18649 15887 18683
rect 15945 18649 15979 18683
rect 16497 18649 16531 18683
rect 17509 18649 17543 18683
rect 3893 18581 3927 18615
rect 8953 18581 8987 18615
rect 16221 18581 16255 18615
rect 19625 18581 19659 18615
rect 26341 18581 26375 18615
rect 4077 18377 4111 18411
rect 9965 18377 9999 18411
rect 13737 18377 13771 18411
rect 15393 18377 15427 18411
rect 15945 18377 15979 18411
rect 16839 18377 16873 18411
rect 17233 18377 17267 18411
rect 18981 18377 19015 18411
rect 19349 18377 19383 18411
rect 2605 18309 2639 18343
rect 16108 18309 16142 18343
rect 16313 18309 16347 18343
rect 17049 18309 17083 18343
rect 19441 18309 19475 18343
rect 2329 18241 2363 18275
rect 10057 18241 10091 18275
rect 13185 18241 13219 18275
rect 14749 18241 14783 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 17325 18241 17359 18275
rect 17601 18241 17635 18275
rect 13461 18173 13495 18207
rect 14381 18173 14415 18207
rect 14657 18173 14691 18207
rect 14841 18173 14875 18207
rect 17509 18173 17543 18207
rect 19533 18173 19567 18207
rect 15117 18105 15151 18139
rect 16681 18105 16715 18139
rect 13553 18037 13587 18071
rect 14749 18037 14783 18071
rect 16129 18037 16163 18071
rect 16865 18037 16899 18071
rect 9965 17833 9999 17867
rect 10333 17833 10367 17867
rect 12725 17833 12759 17867
rect 13461 17833 13495 17867
rect 15485 17833 15519 17867
rect 16957 17833 16991 17867
rect 10701 17765 10735 17799
rect 15025 17697 15059 17731
rect 1409 17629 1443 17663
rect 7021 17629 7055 17663
rect 9689 17629 9723 17663
rect 9781 17629 9815 17663
rect 10057 17629 10091 17663
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 13277 17629 13311 17663
rect 13461 17629 13495 17663
rect 13553 17629 13587 17663
rect 13737 17629 13771 17663
rect 14381 17629 14415 17663
rect 15301 17629 15335 17663
rect 15669 17629 15703 17663
rect 18521 17629 18555 17663
rect 22845 17629 22879 17663
rect 11069 17561 11103 17595
rect 13921 17561 13955 17595
rect 22578 17561 22612 17595
rect 1593 17493 1627 17527
rect 5733 17493 5767 17527
rect 10517 17493 10551 17527
rect 10609 17493 10643 17527
rect 18705 17493 18739 17527
rect 21465 17493 21499 17527
rect 6193 17289 6227 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 12909 17289 12943 17323
rect 15393 17289 15427 17323
rect 18705 17289 18739 17323
rect 9781 17221 9815 17255
rect 13921 17221 13955 17255
rect 14197 17221 14231 17255
rect 18521 17221 18555 17255
rect 20729 17221 20763 17255
rect 3985 17153 4019 17187
rect 4169 17153 4203 17187
rect 4813 17153 4847 17187
rect 5080 17153 5114 17187
rect 6828 17153 6862 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 9873 17153 9907 17187
rect 11529 17153 11563 17187
rect 13185 17153 13219 17187
rect 13461 17153 13495 17187
rect 14841 17153 14875 17187
rect 15945 17153 15979 17187
rect 16865 17153 16899 17187
rect 18797 17153 18831 17187
rect 20821 17153 20855 17187
rect 22845 17153 22879 17187
rect 23029 17153 23063 17187
rect 6561 17085 6595 17119
rect 8493 17085 8527 17119
rect 8861 17085 8895 17119
rect 8953 17085 8987 17119
rect 9689 17085 9723 17119
rect 10885 17085 10919 17119
rect 11161 17085 11195 17119
rect 14657 17085 14691 17119
rect 15669 17085 15703 17119
rect 19073 17085 19107 17119
rect 7941 17017 7975 17051
rect 13553 17017 13587 17051
rect 14473 17017 14507 17051
rect 15025 17017 15059 17051
rect 18153 17017 18187 17051
rect 3985 16949 4019 16983
rect 8401 16949 8435 16983
rect 10241 16949 10275 16983
rect 11713 16949 11747 16983
rect 13093 16949 13127 16983
rect 13921 16949 13955 16983
rect 14105 16949 14139 16983
rect 15761 16949 15795 16983
rect 16773 16949 16807 16983
rect 18521 16949 18555 16983
rect 20545 16949 20579 16983
rect 22845 16949 22879 16983
rect 5273 16745 5307 16779
rect 8769 16745 8803 16779
rect 9781 16745 9815 16779
rect 10425 16745 10459 16779
rect 10977 16745 11011 16779
rect 11621 16745 11655 16779
rect 13461 16745 13495 16779
rect 17049 16745 17083 16779
rect 18521 16745 18555 16779
rect 19441 16745 19475 16779
rect 23121 16745 23155 16779
rect 16865 16677 16899 16711
rect 18889 16677 18923 16711
rect 1685 16609 1719 16643
rect 3801 16609 3835 16643
rect 6285 16609 6319 16643
rect 8217 16609 8251 16643
rect 9505 16609 9539 16643
rect 12449 16609 12483 16643
rect 12817 16609 12851 16643
rect 14105 16609 14139 16643
rect 17141 16609 17175 16643
rect 19533 16609 19567 16643
rect 21649 16609 21683 16643
rect 4068 16541 4102 16575
rect 5273 16541 5307 16575
rect 5457 16541 5491 16575
rect 9873 16541 9907 16575
rect 10149 16541 10183 16575
rect 10701 16541 10735 16575
rect 12357 16541 12391 16575
rect 13093 16541 13127 16575
rect 17417 16541 17451 16575
rect 17509 16541 17543 16575
rect 18337 16541 18371 16575
rect 18613 16541 18647 16575
rect 18705 16541 18739 16575
rect 19257 16541 19291 16575
rect 20453 16541 20487 16575
rect 21557 16541 21591 16575
rect 21741 16541 21775 16575
rect 21833 16541 21867 16575
rect 22569 16541 22603 16575
rect 22753 16541 22787 16575
rect 23673 16541 23707 16575
rect 23857 16541 23891 16575
rect 24041 16541 24075 16575
rect 1952 16473 1986 16507
rect 3341 16473 3375 16507
rect 3525 16473 3559 16507
rect 6552 16473 6586 16507
rect 11253 16473 11287 16507
rect 11437 16473 11471 16507
rect 15025 16473 15059 16507
rect 17693 16473 17727 16507
rect 22937 16473 22971 16507
rect 3065 16405 3099 16439
rect 3157 16405 3191 16439
rect 5181 16405 5215 16439
rect 7665 16405 7699 16439
rect 8953 16405 8987 16439
rect 10609 16405 10643 16439
rect 11161 16405 11195 16439
rect 11897 16405 11931 16439
rect 12265 16405 12299 16439
rect 13001 16405 13035 16439
rect 14749 16405 14783 16439
rect 16313 16405 16347 16439
rect 17877 16405 17911 16439
rect 18061 16405 18095 16439
rect 19809 16405 19843 16439
rect 20361 16405 20395 16439
rect 22477 16405 22511 16439
rect 23949 16405 23983 16439
rect 1593 16201 1627 16235
rect 6837 16201 6871 16235
rect 6929 16201 6963 16235
rect 9873 16201 9907 16235
rect 9965 16201 9999 16235
rect 13829 16201 13863 16235
rect 14289 16201 14323 16235
rect 14381 16201 14415 16235
rect 23949 16201 23983 16235
rect 1930 16133 1964 16167
rect 3893 16133 3927 16167
rect 7097 16133 7131 16167
rect 7297 16133 7331 16167
rect 16849 16133 16883 16167
rect 17049 16133 17083 16167
rect 18705 16133 18739 16167
rect 22100 16133 22134 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 4997 16065 5031 16099
rect 5641 16065 5675 16099
rect 5825 16065 5859 16099
rect 6561 16065 6595 16099
rect 6837 16065 6871 16099
rect 8493 16065 8527 16099
rect 8749 16065 8783 16099
rect 10425 16065 10459 16099
rect 11069 16065 11103 16099
rect 11345 16065 11379 16099
rect 11529 16065 11563 16099
rect 14749 16065 14783 16099
rect 17141 16065 17175 16099
rect 17325 16065 17359 16099
rect 17785 16065 17819 16099
rect 18061 16065 18095 16099
rect 18245 16065 18279 16099
rect 18521 16065 18555 16099
rect 19073 16065 19107 16099
rect 21833 16065 21867 16099
rect 24041 16065 24075 16099
rect 24961 16065 24995 16099
rect 25145 16065 25179 16099
rect 8125 15997 8159 16031
rect 12081 15997 12115 16031
rect 12357 15997 12391 16031
rect 14565 15997 14599 16031
rect 15025 15997 15059 16031
rect 17601 15997 17635 16031
rect 17969 15997 18003 16031
rect 19349 15997 19383 16031
rect 20821 15997 20855 16031
rect 21557 15997 21591 16031
rect 23305 15997 23339 16031
rect 24317 15997 24351 16031
rect 3709 15929 3743 15963
rect 4261 15929 4295 15963
rect 6745 15929 6779 15963
rect 11713 15929 11747 15963
rect 16681 15929 16715 15963
rect 24133 15929 24167 15963
rect 3065 15861 3099 15895
rect 3893 15861 3927 15895
rect 4353 15861 4387 15895
rect 5641 15861 5675 15895
rect 7113 15861 7147 15895
rect 7573 15861 7607 15895
rect 10149 15861 10183 15895
rect 10885 15861 10919 15895
rect 11253 15861 11287 15895
rect 13921 15861 13955 15895
rect 16497 15861 16531 15895
rect 16865 15861 16899 15895
rect 17233 15861 17267 15895
rect 18153 15861 18187 15895
rect 21005 15861 21039 15895
rect 23213 15861 23247 15895
rect 24041 15861 24075 15895
rect 25145 15861 25179 15895
rect 1593 15657 1627 15691
rect 2329 15657 2363 15691
rect 2789 15657 2823 15691
rect 3617 15657 3651 15691
rect 3893 15657 3927 15691
rect 7665 15657 7699 15691
rect 8585 15657 8619 15691
rect 11989 15657 12023 15691
rect 12633 15657 12667 15691
rect 13093 15657 13127 15691
rect 15025 15657 15059 15691
rect 15209 15657 15243 15691
rect 17509 15657 17543 15691
rect 19257 15657 19291 15691
rect 21649 15657 21683 15691
rect 21557 15589 21591 15623
rect 3157 15521 3191 15555
rect 4261 15521 4295 15555
rect 4813 15521 4847 15555
rect 10241 15521 10275 15555
rect 17417 15521 17451 15555
rect 19441 15521 19475 15555
rect 23305 15521 23339 15555
rect 24501 15521 24535 15555
rect 1409 15453 1443 15487
rect 2513 15453 2547 15487
rect 3433 15453 3467 15487
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 5181 15453 5215 15487
rect 7205 15453 7239 15487
rect 7389 15453 7423 15487
rect 7665 15453 7699 15487
rect 7757 15453 7791 15487
rect 8401 15453 8435 15487
rect 8585 15453 8619 15487
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 14933 15453 14967 15487
rect 15117 15453 15151 15487
rect 15669 15453 15703 15487
rect 19533 15453 19567 15487
rect 19901 15453 19935 15487
rect 20729 15453 20763 15487
rect 20821 15453 20855 15487
rect 21649 15453 21683 15487
rect 23049 15453 23083 15487
rect 24041 15453 24075 15487
rect 24768 15453 24802 15487
rect 3249 15385 3283 15419
rect 5448 15385 5482 15419
rect 10517 15385 10551 15419
rect 15393 15385 15427 15419
rect 15577 15385 15611 15419
rect 17693 15385 17727 15419
rect 17877 15385 17911 15419
rect 20085 15385 20119 15419
rect 21373 15385 21407 15419
rect 2605 15317 2639 15351
rect 2789 15317 2823 15351
rect 4445 15317 4479 15351
rect 6561 15317 6595 15351
rect 6653 15317 6687 15351
rect 7481 15317 7515 15351
rect 7849 15317 7883 15351
rect 19625 15317 19659 15351
rect 19809 15317 19843 15351
rect 20913 15317 20947 15351
rect 21925 15317 21959 15351
rect 23397 15317 23431 15351
rect 25881 15317 25915 15351
rect 5641 15113 5675 15147
rect 16681 15113 16715 15147
rect 18061 15113 18095 15147
rect 21005 15113 21039 15147
rect 23765 15113 23799 15147
rect 25145 15113 25179 15147
rect 3065 15045 3099 15079
rect 3281 15045 3315 15079
rect 16221 15045 16255 15079
rect 16405 15045 16439 15079
rect 17877 15045 17911 15079
rect 23397 15045 23431 15079
rect 23613 15045 23647 15079
rect 6009 14977 6043 15011
rect 13093 14977 13127 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 17509 14977 17543 15011
rect 18705 14977 18739 15011
rect 18797 14977 18831 15011
rect 22845 14977 22879 15011
rect 24777 14977 24811 15011
rect 25421 14977 25455 15011
rect 26157 14977 26191 15011
rect 26249 14977 26283 15011
rect 26433 14977 26467 15011
rect 6101 14909 6135 14943
rect 18429 14909 18463 14943
rect 19073 14909 19107 14943
rect 19257 14909 19291 14943
rect 19533 14909 19567 14943
rect 24685 14909 24719 14943
rect 25973 14909 26007 14943
rect 18153 14841 18187 14875
rect 3249 14773 3283 14807
rect 3433 14773 3467 14807
rect 14381 14773 14415 14807
rect 16037 14773 16071 14807
rect 17877 14773 17911 14807
rect 18337 14773 18371 14807
rect 18889 14773 18923 14807
rect 18981 14773 19015 14807
rect 22753 14773 22787 14807
rect 23581 14773 23615 14807
rect 26433 14773 26467 14807
rect 9321 14569 9355 14603
rect 15301 14569 15335 14603
rect 16589 14569 16623 14603
rect 17233 14569 17267 14603
rect 17693 14569 17727 14603
rect 17969 14569 18003 14603
rect 18337 14569 18371 14603
rect 18521 14569 18555 14603
rect 18981 14569 19015 14603
rect 19349 14569 19383 14603
rect 20177 14569 20211 14603
rect 18797 14501 18831 14535
rect 24133 14501 24167 14535
rect 2973 14433 3007 14467
rect 3065 14433 3099 14467
rect 13001 14433 13035 14467
rect 16405 14433 16439 14467
rect 17785 14433 17819 14467
rect 18245 14433 18279 14467
rect 18521 14433 18555 14467
rect 19625 14433 19659 14467
rect 19993 14433 20027 14467
rect 23029 14433 23063 14467
rect 3157 14365 3191 14399
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 4261 14365 4295 14399
rect 4353 14365 4387 14399
rect 4629 14365 4663 14399
rect 6929 14365 6963 14399
rect 7113 14365 7147 14399
rect 7389 14365 7423 14399
rect 7757 14365 7791 14399
rect 7849 14365 7883 14399
rect 8401 14365 8435 14399
rect 8585 14365 8619 14399
rect 9413 14365 9447 14399
rect 9505 14365 9539 14399
rect 9689 14365 9723 14399
rect 14657 14365 14691 14399
rect 14841 14365 14875 14399
rect 15117 14365 15151 14399
rect 15761 14365 15795 14399
rect 16681 14365 16715 14399
rect 16957 14365 16991 14399
rect 17325 14365 17359 14399
rect 17889 14365 17923 14399
rect 18337 14343 18371 14377
rect 18429 14365 18463 14399
rect 19073 14365 19107 14399
rect 19257 14365 19291 14399
rect 19441 14365 19475 14399
rect 22477 14365 22511 14399
rect 22569 14365 22603 14399
rect 22661 14365 22695 14399
rect 22845 14365 22879 14399
rect 23121 14365 23155 14399
rect 23305 14365 23339 14399
rect 23857 14365 23891 14399
rect 24225 14365 24259 14399
rect 24593 14365 24627 14399
rect 4445 14297 4479 14331
rect 8033 14297 8067 14331
rect 12725 14297 12759 14331
rect 15945 14297 15979 14331
rect 23489 14297 23523 14331
rect 23949 14297 23983 14331
rect 24838 14297 24872 14331
rect 2789 14229 2823 14263
rect 3801 14229 3835 14263
rect 4721 14229 4755 14263
rect 7021 14229 7055 14263
rect 7481 14229 7515 14263
rect 8217 14229 8251 14263
rect 8953 14229 8987 14263
rect 9597 14229 9631 14263
rect 12357 14229 12391 14263
rect 12817 14229 12851 14263
rect 14105 14229 14139 14263
rect 14933 14229 14967 14263
rect 15577 14229 15611 14263
rect 16129 14229 16163 14263
rect 16773 14229 16807 14263
rect 17509 14229 17543 14263
rect 19809 14229 19843 14263
rect 22385 14229 22419 14263
rect 23765 14229 23799 14263
rect 24225 14229 24259 14263
rect 25973 14229 26007 14263
rect 1593 14025 1627 14059
rect 3985 14025 4019 14059
rect 6745 14025 6779 14059
rect 7205 14025 7239 14059
rect 8677 14025 8711 14059
rect 9689 14025 9723 14059
rect 13645 14025 13679 14059
rect 14105 14025 14139 14059
rect 14565 14025 14599 14059
rect 15367 14025 15401 14059
rect 18245 14025 18279 14059
rect 22937 14025 22971 14059
rect 24869 14025 24903 14059
rect 26433 14025 26467 14059
rect 2513 13957 2547 13991
rect 6377 13957 6411 13991
rect 7113 13957 7147 13991
rect 10057 13957 10091 13991
rect 14197 13957 14231 13991
rect 15577 13957 15611 13991
rect 22845 13957 22879 13991
rect 23213 13957 23247 13991
rect 25021 13957 25055 13991
rect 25237 13957 25271 13991
rect 6883 13923 6917 13957
rect 1409 13889 1443 13923
rect 2881 13889 2915 13923
rect 4997 13889 5031 13923
rect 5365 13889 5399 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 8125 13889 8159 13923
rect 8309 13889 8343 13923
rect 8401 13889 8435 13923
rect 8493 13889 8527 13923
rect 9781 13889 9815 13923
rect 9873 13889 9907 13923
rect 10793 13889 10827 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 15117 13889 15151 13923
rect 17325 13889 17359 13923
rect 17417 13889 17451 13923
rect 17601 13889 17635 13923
rect 18613 13889 18647 13923
rect 22201 13889 22235 13923
rect 22385 13889 22419 13923
rect 22477 13889 22511 13923
rect 22569 13889 22603 13923
rect 23121 13889 23155 13923
rect 23305 13889 23339 13923
rect 23489 13889 23523 13923
rect 23949 13889 23983 13923
rect 25789 13889 25823 13923
rect 3433 13821 3467 13855
rect 4169 13821 4203 13855
rect 5273 13821 5307 13855
rect 7757 13821 7791 13855
rect 9045 13821 9079 13855
rect 12173 13821 12207 13855
rect 14381 13821 14415 13855
rect 14841 13821 14875 13855
rect 18521 13821 18555 13855
rect 23857 13821 23891 13855
rect 24685 13821 24719 13855
rect 4537 13753 4571 13787
rect 13737 13753 13771 13787
rect 15209 13753 15243 13787
rect 2329 13685 2363 13719
rect 2513 13685 2547 13719
rect 4629 13685 4663 13719
rect 4813 13685 4847 13719
rect 5181 13685 5215 13719
rect 5457 13685 5491 13719
rect 6469 13685 6503 13719
rect 6929 13685 6963 13719
rect 9965 13685 9999 13719
rect 10977 13685 11011 13719
rect 11529 13685 11563 13719
rect 15025 13685 15059 13719
rect 15393 13685 15427 13719
rect 18613 13685 18647 13719
rect 24041 13685 24075 13719
rect 25053 13685 25087 13719
rect 3249 13481 3283 13515
rect 3985 13481 4019 13515
rect 4169 13481 4203 13515
rect 4261 13481 4295 13515
rect 5549 13481 5583 13515
rect 7205 13481 7239 13515
rect 7573 13481 7607 13515
rect 12357 13481 12391 13515
rect 13553 13481 13587 13515
rect 14841 13481 14875 13515
rect 18337 13481 18371 13515
rect 22661 13481 22695 13515
rect 23581 13481 23615 13515
rect 4721 13413 4755 13447
rect 8953 13413 8987 13447
rect 23857 13413 23891 13447
rect 3525 13345 3559 13379
rect 10609 13345 10643 13379
rect 12541 13345 12575 13379
rect 13185 13345 13219 13379
rect 15761 13345 15795 13379
rect 18245 13345 18279 13379
rect 18613 13345 18647 13379
rect 19349 13345 19383 13379
rect 21373 13345 21407 13379
rect 23121 13345 23155 13379
rect 24685 13345 24719 13379
rect 1593 13277 1627 13311
rect 1869 13277 1903 13311
rect 3433 13277 3467 13311
rect 4445 13277 4479 13311
rect 4537 13277 4571 13311
rect 4813 13277 4847 13311
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 5825 13277 5859 13311
rect 6092 13277 6126 13311
rect 7481 13277 7515 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 8401 13277 8435 13311
rect 8493 13277 8527 13311
rect 8585 13277 8619 13311
rect 8769 13277 8803 13311
rect 10066 13277 10100 13311
rect 10333 13277 10367 13311
rect 13645 13277 13679 13311
rect 13921 13277 13955 13311
rect 14841 13277 14875 13311
rect 14933 13277 14967 13311
rect 18337 13277 18371 13311
rect 18705 13277 18739 13311
rect 22845 13277 22879 13311
rect 22937 13277 22971 13311
rect 23213 13277 23247 13311
rect 23765 13277 23799 13311
rect 23949 13277 23983 13311
rect 24041 13277 24075 13311
rect 2114 13209 2148 13243
rect 3801 13209 3835 13243
rect 4001 13209 4035 13243
rect 8033 13209 8067 13243
rect 10885 13209 10919 13243
rect 13829 13209 13863 13243
rect 15853 13209 15887 13243
rect 19625 13209 19659 13243
rect 24952 13209 24986 13243
rect 1777 13141 1811 13175
rect 8125 13141 8159 13175
rect 15209 13141 15243 13175
rect 15945 13141 15979 13175
rect 16313 13141 16347 13175
rect 17969 13141 18003 13175
rect 19073 13141 19107 13175
rect 26065 13141 26099 13175
rect 3249 12937 3283 12971
rect 4905 12937 4939 12971
rect 7757 12937 7791 12971
rect 8033 12937 8067 12971
rect 11529 12937 11563 12971
rect 12541 12937 12575 12971
rect 17969 12937 18003 12971
rect 19809 12937 19843 12971
rect 21005 12937 21039 12971
rect 23765 12937 23799 12971
rect 24317 12937 24351 12971
rect 24869 12937 24903 12971
rect 3985 12869 4019 12903
rect 5273 12869 5307 12903
rect 5365 12869 5399 12903
rect 9321 12869 9355 12903
rect 11069 12869 11103 12903
rect 14749 12869 14783 12903
rect 19993 12869 20027 12903
rect 1869 12801 1903 12835
rect 2136 12801 2170 12835
rect 3433 12801 3467 12835
rect 4445 12801 4479 12835
rect 4721 12801 4755 12835
rect 5181 12801 5215 12835
rect 5549 12801 5583 12835
rect 7665 12801 7699 12835
rect 7941 12801 7975 12835
rect 8217 12801 8251 12835
rect 8401 12801 8435 12835
rect 8677 12801 8711 12835
rect 11345 12801 11379 12835
rect 11897 12801 11931 12835
rect 12725 12801 12759 12835
rect 15209 12801 15243 12835
rect 15669 12801 15703 12835
rect 16129 12801 16163 12835
rect 18061 12801 18095 12835
rect 18889 12801 18923 12835
rect 19717 12801 19751 12835
rect 20913 12801 20947 12835
rect 22017 12801 22051 12835
rect 24777 12801 24811 12835
rect 25053 12801 25087 12835
rect 25329 12801 25363 12835
rect 25513 12801 25547 12835
rect 25789 12801 25823 12835
rect 8493 12733 8527 12767
rect 9597 12733 9631 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 15025 12733 15059 12767
rect 15117 12733 15151 12767
rect 17877 12733 17911 12767
rect 18981 12733 19015 12767
rect 19165 12733 19199 12767
rect 20637 12733 20671 12767
rect 24225 12733 24259 12767
rect 26341 12733 26375 12767
rect 4537 12665 4571 12699
rect 4629 12665 4663 12699
rect 4997 12665 5031 12699
rect 8585 12665 8619 12699
rect 8861 12665 8895 12699
rect 9045 12665 9079 12699
rect 15577 12665 15611 12699
rect 15945 12665 15979 12699
rect 23857 12665 23891 12699
rect 13461 12597 13495 12631
rect 15853 12597 15887 12631
rect 18429 12597 18463 12631
rect 18521 12597 18555 12631
rect 21833 12597 21867 12631
rect 24501 12597 24535 12631
rect 3985 12393 4019 12427
rect 4261 12393 4295 12427
rect 4721 12393 4755 12427
rect 8309 12393 8343 12427
rect 11437 12393 11471 12427
rect 12357 12393 12391 12427
rect 17233 12393 17267 12427
rect 21925 12393 21959 12427
rect 22845 12393 22879 12427
rect 8677 12325 8711 12359
rect 21741 12325 21775 12359
rect 2881 12257 2915 12291
rect 4353 12257 4387 12291
rect 8217 12257 8251 12291
rect 15485 12257 15519 12291
rect 15761 12257 15795 12291
rect 18153 12257 18187 12291
rect 21281 12257 21315 12291
rect 2145 12189 2179 12223
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 3801 12189 3835 12223
rect 4537 12189 4571 12223
rect 8493 12189 8527 12223
rect 11529 12189 11563 12223
rect 13737 12189 13771 12223
rect 17969 12189 18003 12223
rect 18889 12189 18923 12223
rect 19257 12189 19291 12223
rect 23121 12189 23155 12223
rect 13492 12121 13526 12155
rect 19533 12121 19567 12155
rect 21465 12121 21499 12155
rect 17601 12053 17635 12087
rect 18061 12053 18095 12087
rect 18797 12053 18831 12087
rect 22661 12053 22695 12087
rect 14013 11849 14047 11883
rect 16773 11849 16807 11883
rect 17509 11849 17543 11883
rect 20085 11849 20119 11883
rect 16221 11781 16255 11815
rect 17877 11781 17911 11815
rect 19625 11781 19659 11815
rect 22569 11781 22603 11815
rect 24685 11781 24719 11815
rect 13185 11713 13219 11747
rect 16865 11713 16899 11747
rect 17325 11713 17359 11747
rect 19993 11713 20027 11747
rect 21925 11713 21959 11747
rect 22109 11713 22143 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 23213 11713 23247 11747
rect 23397 11713 23431 11747
rect 23673 11713 23707 11747
rect 23949 11713 23983 11747
rect 25237 11713 25271 11747
rect 26525 11713 26559 11747
rect 14105 11645 14139 11679
rect 14289 11645 14323 11679
rect 14473 11645 14507 11679
rect 16497 11645 16531 11679
rect 17601 11645 17635 11679
rect 22937 11645 22971 11679
rect 24777 11645 24811 11679
rect 13645 11577 13679 11611
rect 23489 11577 23523 11611
rect 23765 11577 23799 11611
rect 23857 11577 23891 11611
rect 24225 11577 24259 11611
rect 24317 11577 24351 11611
rect 13001 11509 13035 11543
rect 24961 11509 24995 11543
rect 26341 11509 26375 11543
rect 1593 11305 1627 11339
rect 16129 11305 16163 11339
rect 18705 11305 18739 11339
rect 22017 11305 22051 11339
rect 22937 11305 22971 11339
rect 23673 11305 23707 11339
rect 18337 11237 18371 11271
rect 23489 11237 23523 11271
rect 23857 11237 23891 11271
rect 5181 11169 5215 11203
rect 6929 11169 6963 11203
rect 11805 11169 11839 11203
rect 12081 11169 12115 11203
rect 12357 11169 12391 11203
rect 15945 11169 15979 11203
rect 19257 11169 19291 11203
rect 19533 11169 19567 11203
rect 21281 11169 21315 11203
rect 1409 11101 1443 11135
rect 3249 11101 3283 11135
rect 3525 11101 3559 11135
rect 10149 11101 10183 11135
rect 11529 11101 11563 11135
rect 16037 11101 16071 11135
rect 18153 11101 18187 11135
rect 18521 11101 18555 11135
rect 22109 11101 22143 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 22753 11101 22787 11135
rect 23949 11101 23983 11135
rect 25513 11101 25547 11135
rect 2973 11033 3007 11067
rect 5457 11033 5491 11067
rect 15669 11033 15703 11067
rect 22569 11033 22603 11067
rect 23213 11033 23247 11067
rect 3433 10965 3467 10999
rect 10057 10965 10091 10999
rect 13829 10965 13863 10999
rect 14197 10965 14231 10999
rect 24869 10965 24903 10999
rect 6469 10761 6503 10795
rect 11529 10761 11563 10795
rect 13185 10761 13219 10795
rect 14013 10761 14047 10795
rect 19625 10761 19659 10795
rect 22845 10761 22879 10795
rect 25789 10761 25823 10795
rect 5549 10693 5583 10727
rect 7573 10693 7607 10727
rect 8401 10693 8435 10727
rect 14565 10693 14599 10727
rect 21833 10693 21867 10727
rect 22445 10693 22479 10727
rect 22661 10693 22695 10727
rect 24317 10693 24351 10727
rect 24654 10693 24688 10727
rect 1593 10625 1627 10659
rect 3893 10625 3927 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 4353 10625 4387 10659
rect 4813 10625 4847 10659
rect 4997 10625 5031 10659
rect 5089 10625 5123 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 6561 10625 6595 10659
rect 7389 10625 7423 10659
rect 8125 10625 8159 10659
rect 8493 10625 8527 10659
rect 8677 10625 8711 10659
rect 11345 10625 11379 10659
rect 13093 10625 13127 10659
rect 13829 10625 13863 10659
rect 15025 10625 15059 10659
rect 19533 10625 19567 10659
rect 22017 10625 22051 10659
rect 22937 10625 22971 10659
rect 23857 10625 23891 10659
rect 24133 10625 24167 10659
rect 24409 10625 24443 10659
rect 1869 10557 1903 10591
rect 3617 10557 3651 10591
rect 8309 10557 8343 10591
rect 9045 10557 9079 10591
rect 9321 10557 9355 10591
rect 11069 10557 11103 10591
rect 12081 10557 12115 10591
rect 14657 10557 14691 10591
rect 14749 10557 14783 10591
rect 15209 10557 15243 10591
rect 4169 10489 4203 10523
rect 4537 10489 4571 10523
rect 5365 10489 5399 10523
rect 7941 10489 7975 10523
rect 14197 10489 14231 10523
rect 3801 10421 3835 10455
rect 4629 10421 4663 10455
rect 5181 10421 5215 10455
rect 7757 10421 7791 10455
rect 8401 10421 8435 10455
rect 8493 10421 8527 10455
rect 11253 10421 11287 10455
rect 22201 10421 22235 10455
rect 22293 10421 22327 10455
rect 22477 10421 22511 10455
rect 23949 10421 23983 10455
rect 5549 10217 5583 10251
rect 5641 10217 5675 10251
rect 8309 10217 8343 10251
rect 11437 10217 11471 10251
rect 14565 10217 14599 10251
rect 22293 10217 22327 10251
rect 9275 10149 9309 10183
rect 13737 10149 13771 10183
rect 14381 10149 14415 10183
rect 22017 10149 22051 10183
rect 1593 10081 1627 10115
rect 5089 10081 5123 10115
rect 7389 10081 7423 10115
rect 7665 10081 7699 10115
rect 9689 10081 9723 10115
rect 11621 10081 11655 10115
rect 22753 10081 22787 10115
rect 24685 10081 24719 10115
rect 4169 10013 4203 10047
rect 4629 10013 4663 10047
rect 4905 10013 4939 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 6101 10013 6135 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7297 10013 7331 10047
rect 7757 10013 7791 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 13553 10013 13587 10047
rect 14197 10013 14231 10047
rect 14473 10013 14507 10047
rect 20637 10013 20671 10047
rect 22661 10013 22695 10047
rect 22937 10013 22971 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 26341 10013 26375 10047
rect 1869 9945 1903 9979
rect 3617 9945 3651 9979
rect 4261 9945 4295 9979
rect 4353 9945 4387 9979
rect 4491 9945 4525 9979
rect 4721 9945 4755 9979
rect 5825 9945 5859 9979
rect 6469 9945 6503 9979
rect 8033 9945 8067 9979
rect 9045 9945 9079 9979
rect 9965 9945 9999 9979
rect 11897 9945 11931 9979
rect 20904 9945 20938 9979
rect 22293 9945 22327 9979
rect 24952 9945 24986 9979
rect 3985 9877 4019 9911
rect 6653 9877 6687 9911
rect 7021 9877 7055 9911
rect 8401 9877 8435 9911
rect 13369 9877 13403 9911
rect 22109 9877 22143 9911
rect 23121 9877 23155 9911
rect 24593 9877 24627 9911
rect 26065 9877 26099 9911
rect 26157 9877 26191 9911
rect 4997 9673 5031 9707
rect 5825 9673 5859 9707
rect 21281 9673 21315 9707
rect 21925 9673 21959 9707
rect 24041 9673 24075 9707
rect 25329 9673 25363 9707
rect 5977 9605 6011 9639
rect 6193 9605 6227 9639
rect 6745 9605 6779 9639
rect 7849 9605 7883 9639
rect 7941 9605 7975 9639
rect 10241 9605 10275 9639
rect 11621 9605 11655 9639
rect 22385 9605 22419 9639
rect 23673 9605 23707 9639
rect 23889 9605 23923 9639
rect 24961 9605 24995 9639
rect 25177 9605 25211 9639
rect 25789 9605 25823 9639
rect 6515 9571 6549 9605
rect 2329 9537 2363 9571
rect 4445 9537 4479 9571
rect 4721 9537 4755 9571
rect 5549 9537 5583 9571
rect 7021 9537 7055 9571
rect 7665 9537 7699 9571
rect 8033 9537 8067 9571
rect 8493 9537 8527 9571
rect 8585 9537 8619 9571
rect 8677 9537 8711 9571
rect 8769 9537 8803 9571
rect 10333 9537 10367 9571
rect 11529 9537 11563 9571
rect 14657 9537 14691 9571
rect 18521 9537 18555 9571
rect 21465 9537 21499 9571
rect 22109 9537 22143 9571
rect 22569 9537 22603 9571
rect 23029 9537 23063 9571
rect 23305 9537 23339 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 2697 9469 2731 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 4629 9469 4663 9503
rect 5273 9469 5307 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 8309 9469 8343 9503
rect 15025 9469 15059 9503
rect 18153 9469 18187 9503
rect 22753 9469 22787 9503
rect 22845 9469 22879 9503
rect 22937 9469 22971 9503
rect 23489 9401 23523 9435
rect 4123 9333 4157 9367
rect 5457 9333 5491 9367
rect 6009 9333 6043 9367
rect 6377 9333 6411 9367
rect 6561 9333 6595 9367
rect 8217 9333 8251 9367
rect 16451 9333 16485 9367
rect 16773 9333 16807 9367
rect 22201 9333 22235 9367
rect 23213 9333 23247 9367
rect 23857 9333 23891 9367
rect 25145 9333 25179 9367
rect 2789 9129 2823 9163
rect 6009 9129 6043 9163
rect 7481 9129 7515 9163
rect 10977 9129 11011 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 13461 9129 13495 9163
rect 15669 9129 15703 9163
rect 16681 9129 16715 9163
rect 17509 9129 17543 9163
rect 18889 9129 18923 9163
rect 21741 9129 21775 9163
rect 23673 9129 23707 9163
rect 4353 9061 4387 9095
rect 12357 9061 12391 9095
rect 17417 9061 17451 9095
rect 23489 9061 23523 9095
rect 24041 9061 24075 9095
rect 4077 8993 4111 9027
rect 7849 8993 7883 9027
rect 17141 8993 17175 9027
rect 18153 8993 18187 9027
rect 18245 8993 18279 9027
rect 22017 8993 22051 9027
rect 1409 8925 1443 8959
rect 2881 8925 2915 8959
rect 3985 8925 4019 8959
rect 6101 8925 6135 8959
rect 7665 8925 7699 8959
rect 15577 8925 15611 8959
rect 16589 8925 16623 8959
rect 17049 8925 17083 8959
rect 17693 8925 17727 8959
rect 17877 8925 17911 8959
rect 19441 8925 19475 8959
rect 20637 8925 20671 8959
rect 21373 8925 21407 8959
rect 25789 8925 25823 8959
rect 10793 8857 10827 8891
rect 12509 8857 12543 8891
rect 12725 8857 12759 8891
rect 12969 8857 13003 8891
rect 13185 8857 13219 8891
rect 13277 8857 13311 8891
rect 13477 8857 13511 8891
rect 17785 8857 17819 8891
rect 18015 8857 18049 8891
rect 18429 8857 18463 8891
rect 18613 8857 18647 8891
rect 18705 8857 18739 8891
rect 18910 8857 18944 8891
rect 22284 8857 22318 8891
rect 1593 8789 1627 8823
rect 10993 8789 11027 8823
rect 11161 8789 11195 8823
rect 12817 8789 12851 8823
rect 13645 8789 13679 8823
rect 19073 8789 19107 8823
rect 19349 8789 19383 8823
rect 20545 8789 20579 8823
rect 21741 8789 21775 8823
rect 21925 8789 21959 8823
rect 23397 8789 23431 8823
rect 23673 8789 23707 8823
rect 25697 8789 25731 8823
rect 8743 8585 8777 8619
rect 13645 8585 13679 8619
rect 17141 8585 17175 8619
rect 18429 8585 18463 8619
rect 22477 8585 22511 8619
rect 22753 8585 22787 8619
rect 8953 8517 8987 8551
rect 13369 8517 13403 8551
rect 14105 8517 14139 8551
rect 23866 8517 23900 8551
rect 13093 8449 13127 8483
rect 14013 8449 14047 8483
rect 15209 8449 15243 8483
rect 17969 8449 18003 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 18889 8449 18923 8483
rect 19165 8449 19199 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 22661 8449 22695 8483
rect 24133 8449 24167 8483
rect 13277 8381 13311 8415
rect 15393 8381 15427 8415
rect 17325 8381 17359 8415
rect 17417 8381 17451 8415
rect 17509 8381 17543 8415
rect 17601 8381 17635 8415
rect 17785 8381 17819 8415
rect 18153 8381 18187 8415
rect 18797 8381 18831 8415
rect 19809 8381 19843 8415
rect 8585 8313 8619 8347
rect 12909 8313 12943 8347
rect 13461 8313 13495 8347
rect 14381 8313 14415 8347
rect 18061 8313 18095 8347
rect 18705 8313 18739 8347
rect 8769 8245 8803 8279
rect 13369 8245 13403 8279
rect 13645 8245 13679 8279
rect 14565 8245 14599 8279
rect 21235 8245 21269 8279
rect 5549 8041 5583 8075
rect 12081 8041 12115 8075
rect 12817 8041 12851 8075
rect 13369 8041 13403 8075
rect 13553 8041 13587 8075
rect 14105 8041 14139 8075
rect 18153 8041 18187 8075
rect 18337 8041 18371 8075
rect 19809 8041 19843 8075
rect 11069 7973 11103 8007
rect 12633 7973 12667 8007
rect 14473 7973 14507 8007
rect 2237 7905 2271 7939
rect 4077 7905 4111 7939
rect 12265 7905 12299 7939
rect 13185 7905 13219 7939
rect 13921 7905 13955 7939
rect 18429 7905 18463 7939
rect 18889 7905 18923 7939
rect 19993 7905 20027 7939
rect 20085 7905 20119 7939
rect 20177 7905 20211 7939
rect 2145 7837 2179 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 7941 7837 7975 7871
rect 9137 7837 9171 7871
rect 11345 7837 11379 7871
rect 11437 7837 11471 7871
rect 11621 7837 11655 7871
rect 12081 7837 12115 7871
rect 12357 7837 12391 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14652 7837 14686 7871
rect 15024 7837 15058 7871
rect 15117 7837 15151 7871
rect 15347 7837 15381 7871
rect 15760 7837 15794 7871
rect 15853 7837 15887 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 18981 7837 19015 7871
rect 19257 7837 19291 7871
rect 19533 7837 19567 7871
rect 19625 7837 19659 7871
rect 20269 7837 20303 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 7757 7769 7791 7803
rect 7849 7769 7883 7803
rect 8953 7769 8987 7803
rect 9321 7769 9355 7803
rect 11069 7769 11103 7803
rect 11253 7769 11287 7803
rect 13553 7769 13587 7803
rect 14749 7769 14783 7803
rect 14841 7769 14875 7803
rect 15485 7769 15519 7803
rect 15577 7769 15611 7803
rect 19441 7769 19475 7803
rect 3893 7701 3927 7735
rect 8125 7701 8159 7735
rect 11529 7701 11563 7735
rect 12541 7701 12575 7735
rect 12817 7701 12851 7735
rect 15209 7701 15243 7735
rect 20453 7701 20487 7735
rect 20913 7701 20947 7735
rect 4537 7497 4571 7531
rect 7481 7497 7515 7531
rect 7941 7497 7975 7531
rect 11897 7497 11931 7531
rect 11989 7497 12023 7531
rect 13369 7497 13403 7531
rect 14749 7497 14783 7531
rect 17233 7497 17267 7531
rect 17877 7497 17911 7531
rect 19533 7497 19567 7531
rect 21189 7497 21223 7531
rect 21281 7497 21315 7531
rect 5641 7429 5675 7463
rect 8493 7429 8527 7463
rect 8769 7429 8803 7463
rect 12173 7429 12207 7463
rect 13829 7429 13863 7463
rect 14289 7429 14323 7463
rect 20269 7429 20303 7463
rect 21433 7429 21467 7463
rect 21649 7429 21683 7463
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4997 7361 5031 7395
rect 5457 7361 5491 7395
rect 5733 7361 5767 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 7849 7361 7883 7395
rect 8309 7361 8343 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 9137 7361 9171 7395
rect 9689 7361 9723 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 13001 7361 13035 7395
rect 16773 7361 16807 7395
rect 17049 7361 17083 7395
rect 17417 7361 17451 7395
rect 17877 7361 17911 7395
rect 18245 7361 18279 7395
rect 20085 7361 20119 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 20821 7361 20855 7395
rect 21005 7361 21039 7395
rect 5089 7293 5123 7327
rect 8125 7293 8159 7327
rect 9229 7293 9263 7327
rect 9505 7293 9539 7327
rect 10149 7293 10183 7327
rect 10425 7293 10459 7327
rect 10563 7293 10597 7327
rect 10701 7293 10735 7327
rect 16865 7293 16899 7327
rect 12541 7225 12575 7259
rect 14197 7225 14231 7259
rect 14565 7225 14599 7259
rect 17693 7225 17727 7259
rect 3065 7157 3099 7191
rect 4721 7157 4755 7191
rect 5273 7157 5307 7191
rect 5825 7157 5859 7191
rect 7389 7157 7423 7191
rect 9413 7157 9447 7191
rect 11345 7157 11379 7191
rect 12173 7157 12207 7191
rect 13369 7157 13403 7191
rect 13553 7157 13587 7191
rect 13645 7157 13679 7191
rect 13829 7157 13863 7191
rect 16773 7157 16807 7191
rect 17555 7157 17589 7191
rect 20637 7157 20671 7191
rect 21465 7157 21499 7191
rect 5273 6953 5307 6987
rect 8217 6953 8251 6987
rect 8677 6953 8711 6987
rect 9045 6953 9079 6987
rect 9505 6953 9539 6987
rect 10333 6953 10367 6987
rect 10793 6953 10827 6987
rect 11621 6953 11655 6987
rect 12357 6953 12391 6987
rect 13645 6953 13679 6987
rect 20545 6953 20579 6987
rect 10241 6885 10275 6919
rect 1593 6817 1627 6851
rect 3341 6817 3375 6851
rect 4077 6817 4111 6851
rect 4721 6817 4755 6851
rect 5733 6817 5767 6851
rect 5825 6817 5859 6851
rect 9229 6817 9263 6851
rect 9965 6817 9999 6851
rect 13645 6817 13679 6851
rect 15853 6817 15887 6851
rect 19073 6817 19107 6851
rect 20269 6817 20303 6851
rect 21005 6817 21039 6851
rect 22477 6817 22511 6851
rect 3617 6749 3651 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 5641 6749 5675 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 8953 6749 8987 6783
rect 9781 6749 9815 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 10517 6749 10551 6783
rect 10609 6749 10643 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 11805 6749 11839 6783
rect 12081 6749 12115 6783
rect 13553 6749 13587 6783
rect 13829 6749 13863 6783
rect 16221 6749 16255 6783
rect 17647 6749 17681 6783
rect 18337 6749 18371 6783
rect 18705 6749 18739 6783
rect 18889 6749 18923 6783
rect 19257 6749 19291 6783
rect 19901 6749 19935 6783
rect 20177 6749 20211 6783
rect 20637 6749 20671 6783
rect 4353 6681 4387 6715
rect 4445 6681 4479 6715
rect 4583 6681 4617 6715
rect 5457 6681 5491 6715
rect 10977 6681 11011 6715
rect 12341 6681 12375 6715
rect 12541 6681 12575 6715
rect 17785 6681 17819 6715
rect 3893 6613 3927 6647
rect 4813 6613 4847 6647
rect 6101 6613 6135 6647
rect 11989 6613 12023 6647
rect 12173 6613 12207 6647
rect 13369 6613 13403 6647
rect 1593 6409 1627 6443
rect 2421 6409 2455 6443
rect 4445 6409 4479 6443
rect 7113 6409 7147 6443
rect 8033 6409 8067 6443
rect 9337 6409 9371 6443
rect 10349 6409 10383 6443
rect 10701 6409 10735 6443
rect 16313 6409 16347 6443
rect 16957 6409 16991 6443
rect 20637 6409 20671 6443
rect 21925 6409 21959 6443
rect 5549 6341 5583 6375
rect 5825 6341 5859 6375
rect 5917 6341 5951 6375
rect 7573 6341 7607 6375
rect 7665 6341 7699 6375
rect 8125 6341 8159 6375
rect 8585 6341 8619 6375
rect 9137 6341 9171 6375
rect 9597 6341 9631 6375
rect 10149 6341 10183 6375
rect 19901 6341 19935 6375
rect 1409 6273 1443 6307
rect 2145 6273 2179 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 4905 6273 4939 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 5641 6273 5675 6307
rect 6009 6273 6043 6307
rect 6745 6273 6779 6307
rect 7297 6273 7331 6307
rect 7849 6273 7883 6307
rect 8309 6273 8343 6307
rect 8493 6273 8527 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9873 6273 9907 6307
rect 10609 6273 10643 6307
rect 10793 6273 10827 6307
rect 15209 6273 15243 6307
rect 16405 6273 16439 6307
rect 17049 6273 17083 6307
rect 19257 6273 19291 6307
rect 19441 6273 19475 6307
rect 19717 6273 19751 6307
rect 20821 6273 20855 6307
rect 21281 6273 21315 6307
rect 21833 6273 21867 6307
rect 3893 6205 3927 6239
rect 4721 6205 4755 6239
rect 6377 6205 6411 6239
rect 6561 6205 6595 6239
rect 6653 6205 6687 6239
rect 6837 6205 6871 6239
rect 7481 6205 7515 6239
rect 9781 6205 9815 6239
rect 19349 6205 19383 6239
rect 21189 6205 21223 6239
rect 9505 6137 9539 6171
rect 10517 6137 10551 6171
rect 20913 6137 20947 6171
rect 2237 6069 2271 6103
rect 6193 6069 6227 6103
rect 7297 6069 7331 6103
rect 9321 6069 9355 6103
rect 9873 6069 9907 6103
rect 10057 6069 10091 6103
rect 10333 6069 10367 6103
rect 15117 6069 15151 6103
rect 19533 6069 19567 6103
rect 5181 5865 5215 5899
rect 5549 5865 5583 5899
rect 6193 5865 6227 5899
rect 9689 5865 9723 5899
rect 25697 5865 25731 5899
rect 4997 5797 5031 5831
rect 6423 5797 6457 5831
rect 9597 5797 9631 5831
rect 14151 5797 14185 5831
rect 19349 5797 19383 5831
rect 5641 5661 5675 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 6561 5661 6595 5695
rect 9321 5661 9355 5695
rect 9413 5661 9447 5695
rect 9965 5661 9999 5695
rect 15577 5661 15611 5695
rect 15945 5661 15979 5695
rect 19349 5661 19383 5695
rect 19533 5661 19567 5695
rect 19625 5661 19659 5695
rect 19717 5661 19751 5695
rect 19901 5661 19935 5695
rect 25789 5661 25823 5695
rect 5165 5593 5199 5627
rect 5365 5593 5399 5627
rect 9597 5593 9631 5627
rect 9689 5593 9723 5627
rect 9873 5593 9907 5627
rect 16037 5593 16071 5627
rect 17785 5593 17819 5627
rect 19809 5593 19843 5627
rect 5825 5321 5859 5355
rect 5993 5321 6027 5355
rect 14289 5321 14323 5355
rect 6193 5253 6227 5287
rect 9597 5253 9631 5287
rect 13645 5253 13679 5287
rect 19165 5253 19199 5287
rect 2145 5185 2179 5219
rect 2421 5185 2455 5219
rect 2513 5185 2547 5219
rect 12449 5185 12483 5219
rect 12633 5185 12667 5219
rect 13277 5185 13311 5219
rect 13553 5185 13587 5219
rect 13737 5185 13771 5219
rect 13829 5185 13863 5219
rect 14105 5185 14139 5219
rect 14657 5185 14691 5219
rect 15117 5185 15151 5219
rect 15301 5185 15335 5219
rect 19349 5185 19383 5219
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 2237 5117 2271 5151
rect 13921 5117 13955 5151
rect 14565 5117 14599 5151
rect 14749 5117 14783 5151
rect 14841 5117 14875 5151
rect 13415 5049 13449 5083
rect 6009 4981 6043 5015
rect 8309 4981 8343 5015
rect 12633 4981 12667 5015
rect 14105 4981 14139 5015
rect 15025 4981 15059 5015
rect 15209 4981 15243 5015
rect 19165 4981 19199 5015
rect 19993 4981 20027 5015
rect 1593 4777 1627 4811
rect 8125 4777 8159 4811
rect 13737 4777 13771 4811
rect 14657 4777 14691 4811
rect 16497 4777 16531 4811
rect 21051 4777 21085 4811
rect 6653 4641 6687 4675
rect 10149 4641 10183 4675
rect 10517 4641 10551 4675
rect 14749 4641 14783 4675
rect 16313 4641 16347 4675
rect 16957 4641 16991 4675
rect 17049 4641 17083 4675
rect 17141 4641 17175 4675
rect 19257 4641 19291 4675
rect 19625 4641 19659 4675
rect 1409 4573 1443 4607
rect 4813 4573 4847 4607
rect 4997 4573 5031 4607
rect 6377 4573 6411 4607
rect 8401 4573 8435 4607
rect 10057 4573 10091 4607
rect 11943 4573 11977 4607
rect 12725 4573 12759 4607
rect 13001 4573 13035 4607
rect 13093 4573 13127 4607
rect 13277 4573 13311 4607
rect 13461 4573 13495 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 14933 4573 14967 4607
rect 15209 4573 15243 4607
rect 15853 4573 15887 4607
rect 16221 4573 16255 4607
rect 16865 4573 16899 4607
rect 17509 4573 17543 4607
rect 5365 4505 5399 4539
rect 5549 4505 5583 4539
rect 5733 4505 5767 4539
rect 8309 4505 8343 4539
rect 12817 4505 12851 4539
rect 13553 4505 13587 4539
rect 14381 4505 14415 4539
rect 18061 4505 18095 4539
rect 18245 4505 18279 4539
rect 4905 4437 4939 4471
rect 9965 4437 9999 4471
rect 12541 4437 12575 4471
rect 13369 4437 13403 4471
rect 13753 4437 13787 4471
rect 13921 4437 13955 4471
rect 15117 4437 15151 4471
rect 15761 4437 15795 4471
rect 16681 4437 16715 4471
rect 17417 4437 17451 4471
rect 18429 4437 18463 4471
rect 4261 4233 4295 4267
rect 10609 4233 10643 4267
rect 11982 4233 12016 4267
rect 14999 4233 15033 4267
rect 18153 4233 18187 4267
rect 20591 4233 20625 4267
rect 4077 4165 4111 4199
rect 4721 4165 4755 4199
rect 5089 4165 5123 4199
rect 6009 4165 6043 4199
rect 10241 4165 10275 4199
rect 12081 4165 12115 4199
rect 12357 4165 12391 4199
rect 13461 4165 13495 4199
rect 15209 4165 15243 4199
rect 16773 4165 16807 4199
rect 17692 4165 17726 4199
rect 20821 4165 20855 4199
rect 4353 4097 4387 4131
rect 4445 4097 4479 4131
rect 4537 4097 4571 4131
rect 4997 4097 5031 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 6561 4097 6595 4131
rect 6745 4097 6779 4131
rect 8125 4097 8159 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 11529 4097 11563 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 12541 4097 12575 4131
rect 12817 4097 12851 4131
rect 13277 4097 13311 4131
rect 15301 4097 15335 4131
rect 15669 4097 15703 4131
rect 16957 4097 16991 4131
rect 17049 4097 17083 4131
rect 17233 4097 17267 4131
rect 17575 4097 17609 4131
rect 17785 4097 17819 4131
rect 17877 4097 17911 4131
rect 18337 4097 18371 4131
rect 18429 4097 18463 4131
rect 18613 4097 18647 4131
rect 18797 4097 18831 4131
rect 19165 4097 19199 4131
rect 20913 4097 20947 4131
rect 26525 4097 26559 4131
rect 8401 4029 8435 4063
rect 10149 4029 10183 4063
rect 11161 4029 11195 4063
rect 12173 4029 12207 4063
rect 12909 4029 12943 4063
rect 13185 4029 13219 4063
rect 17417 4029 17451 4063
rect 18521 4029 18555 4063
rect 4905 3961 4939 3995
rect 14841 3961 14875 3995
rect 15853 3961 15887 3995
rect 17141 3961 17175 3995
rect 26341 3961 26375 3995
rect 4077 3893 4111 3927
rect 4721 3893 4755 3927
rect 6193 3893 6227 3927
rect 6377 3893 6411 3927
rect 10241 3893 10275 3927
rect 11621 3893 11655 3927
rect 13645 3893 13679 3927
rect 15025 3893 15059 3927
rect 15485 3893 15519 3927
rect 18061 3893 18095 3927
rect 5549 3689 5583 3723
rect 9045 3689 9079 3723
rect 11851 3689 11885 3723
rect 14197 3689 14231 3723
rect 16313 3689 16347 3723
rect 13737 3621 13771 3655
rect 3801 3553 3835 3587
rect 6745 3553 6779 3587
rect 10057 3553 10091 3587
rect 10425 3553 10459 3587
rect 12817 3553 12851 3587
rect 13093 3553 13127 3587
rect 15577 3553 15611 3587
rect 15945 3553 15979 3587
rect 18061 3553 18095 3587
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 5825 3485 5859 3519
rect 8953 3485 8987 3519
rect 9781 3485 9815 3519
rect 12725 3485 12759 3519
rect 13185 3485 13219 3519
rect 13369 3485 13403 3519
rect 13553 3485 13587 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 18613 3485 18647 3519
rect 7021 3417 7055 3451
rect 8769 3417 8803 3451
rect 13461 3417 13495 3451
rect 3525 3349 3559 3383
rect 6469 3349 6503 3383
rect 9229 3349 9263 3383
rect 18245 3349 18279 3383
rect 18521 3349 18555 3383
rect 6929 3145 6963 3179
rect 7941 3145 7975 3179
rect 8493 3145 8527 3179
rect 8861 3145 8895 3179
rect 10839 3145 10873 3179
rect 14841 3145 14875 3179
rect 18429 3145 18463 3179
rect 6561 3077 6595 3111
rect 16957 3077 16991 3111
rect 3709 3009 3743 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 8585 3009 8619 3043
rect 8769 3009 8803 3043
rect 14933 3009 14967 3043
rect 16681 3009 16715 3043
rect 3985 2941 4019 2975
rect 5641 2941 5675 2975
rect 6101 2941 6135 2975
rect 7021 2941 7055 2975
rect 7297 2941 7331 2975
rect 9045 2941 9079 2975
rect 9413 2941 9447 2975
rect 5457 2805 5491 2839
rect 1593 2601 1627 2635
rect 5733 2601 5767 2635
rect 9597 2601 9631 2635
rect 1409 2397 1443 2431
rect 5733 2397 5767 2431
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 9505 2397 9539 2431
rect 10425 2397 10459 2431
rect 14473 2397 14507 2431
rect 18061 2397 18095 2431
rect 25973 2397 26007 2431
rect 6377 2329 6411 2363
rect 10057 2329 10091 2363
rect 14105 2329 14139 2363
rect 22017 2329 22051 2363
rect 18153 2261 18187 2295
rect 22109 2261 22143 2295
rect 26065 2261 26099 2295
<< metal1 >>
rect 1104 27770 26864 27792
rect 1104 27718 4169 27770
rect 4221 27718 4233 27770
rect 4285 27718 4297 27770
rect 4349 27718 4361 27770
rect 4413 27718 4425 27770
rect 4477 27718 10608 27770
rect 10660 27718 10672 27770
rect 10724 27718 10736 27770
rect 10788 27718 10800 27770
rect 10852 27718 10864 27770
rect 10916 27718 17047 27770
rect 17099 27718 17111 27770
rect 17163 27718 17175 27770
rect 17227 27718 17239 27770
rect 17291 27718 17303 27770
rect 17355 27718 23486 27770
rect 23538 27718 23550 27770
rect 23602 27718 23614 27770
rect 23666 27718 23678 27770
rect 23730 27718 23742 27770
rect 23794 27718 26864 27770
rect 1104 27696 26864 27718
rect 3418 27548 3424 27600
rect 3476 27588 3482 27600
rect 3881 27591 3939 27597
rect 3881 27588 3893 27591
rect 3476 27560 3893 27588
rect 3476 27548 3482 27560
rect 3881 27557 3893 27560
rect 3927 27557 3939 27591
rect 3881 27551 3939 27557
rect 10410 27548 10416 27600
rect 10468 27588 10474 27600
rect 10597 27591 10655 27597
rect 10597 27588 10609 27591
rect 10468 27560 10609 27588
rect 10468 27548 10474 27560
rect 10597 27557 10609 27560
rect 10643 27557 10655 27591
rect 10597 27551 10655 27557
rect 17402 27548 17408 27600
rect 17460 27588 17466 27600
rect 17773 27591 17831 27597
rect 17773 27588 17785 27591
rect 17460 27560 17785 27588
rect 17460 27548 17466 27560
rect 17773 27557 17785 27560
rect 17819 27557 17831 27591
rect 17773 27551 17831 27557
rect 24854 27548 24860 27600
rect 24912 27548 24918 27600
rect 4157 27387 4215 27393
rect 4157 27353 4169 27387
rect 4203 27384 4215 27387
rect 5350 27384 5356 27396
rect 4203 27356 5356 27384
rect 4203 27353 4215 27356
rect 4157 27347 4215 27353
rect 5350 27344 5356 27356
rect 5408 27344 5414 27396
rect 6917 27387 6975 27393
rect 6917 27353 6929 27387
rect 6963 27384 6975 27387
rect 7006 27384 7012 27396
rect 6963 27356 7012 27384
rect 6963 27353 6975 27356
rect 6917 27347 6975 27353
rect 7006 27344 7012 27356
rect 7064 27344 7070 27396
rect 7098 27344 7104 27396
rect 7156 27344 7162 27396
rect 10410 27344 10416 27396
rect 10468 27384 10474 27396
rect 10873 27387 10931 27393
rect 10873 27384 10885 27387
rect 10468 27356 10885 27384
rect 10468 27344 10474 27356
rect 10873 27353 10885 27356
rect 10919 27353 10931 27387
rect 10873 27347 10931 27353
rect 16574 27344 16580 27396
rect 16632 27384 16638 27396
rect 17589 27387 17647 27393
rect 17589 27384 17601 27387
rect 16632 27356 17601 27384
rect 16632 27344 16638 27356
rect 17589 27353 17601 27356
rect 17635 27353 17647 27387
rect 17589 27347 17647 27353
rect 24578 27344 24584 27396
rect 24636 27344 24642 27396
rect 4338 27276 4344 27328
rect 4396 27316 4402 27328
rect 6733 27319 6791 27325
rect 6733 27316 6745 27319
rect 4396 27288 6745 27316
rect 4396 27276 4402 27288
rect 6733 27285 6745 27288
rect 6779 27285 6791 27319
rect 6733 27279 6791 27285
rect 1104 27226 26864 27248
rect 1104 27174 4829 27226
rect 4881 27174 4893 27226
rect 4945 27174 4957 27226
rect 5009 27174 5021 27226
rect 5073 27174 5085 27226
rect 5137 27174 11268 27226
rect 11320 27174 11332 27226
rect 11384 27174 11396 27226
rect 11448 27174 11460 27226
rect 11512 27174 11524 27226
rect 11576 27174 17707 27226
rect 17759 27174 17771 27226
rect 17823 27174 17835 27226
rect 17887 27174 17899 27226
rect 17951 27174 17963 27226
rect 18015 27174 24146 27226
rect 24198 27174 24210 27226
rect 24262 27174 24274 27226
rect 24326 27174 24338 27226
rect 24390 27174 24402 27226
rect 24454 27174 26864 27226
rect 1104 27152 26864 27174
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 4249 27115 4307 27121
rect 4249 27112 4261 27115
rect 4212 27084 4261 27112
rect 4212 27072 4218 27084
rect 4249 27081 4261 27084
rect 4295 27112 4307 27115
rect 14826 27112 14832 27124
rect 4295 27084 6684 27112
rect 4295 27081 4307 27084
rect 4249 27075 4307 27081
rect 4338 27044 4344 27056
rect 4172 27016 4344 27044
rect 3326 26936 3332 26988
rect 3384 26976 3390 26988
rect 4172 26985 4200 27016
rect 4338 27004 4344 27016
rect 4396 27004 4402 27056
rect 4157 26979 4215 26985
rect 4157 26976 4169 26979
rect 3384 26948 4169 26976
rect 3384 26936 3390 26948
rect 4157 26945 4169 26948
rect 4203 26945 4215 26979
rect 4157 26939 4215 26945
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26976 4491 26979
rect 4525 26979 4583 26985
rect 4525 26976 4537 26979
rect 4479 26948 4537 26976
rect 4479 26945 4491 26948
rect 4433 26939 4491 26945
rect 4525 26945 4537 26948
rect 4571 26976 4583 26979
rect 6362 26976 6368 26988
rect 4571 26948 6368 26976
rect 4571 26945 4583 26948
rect 4525 26939 4583 26945
rect 6362 26936 6368 26948
rect 6420 26976 6426 26988
rect 6549 26979 6607 26985
rect 6549 26976 6561 26979
rect 6420 26948 6561 26976
rect 6420 26936 6426 26948
rect 6549 26945 6561 26948
rect 6595 26945 6607 26979
rect 6656 26976 6684 27084
rect 10980 27084 14832 27112
rect 6733 27047 6791 27053
rect 6733 27013 6745 27047
rect 6779 27044 6791 27047
rect 7561 27047 7619 27053
rect 7561 27044 7573 27047
rect 6779 27016 7573 27044
rect 6779 27013 6791 27016
rect 6733 27007 6791 27013
rect 7561 27013 7573 27016
rect 7607 27013 7619 27047
rect 7561 27007 7619 27013
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 6656 26948 6837 26976
rect 6549 26939 6607 26945
rect 6825 26945 6837 26948
rect 6871 26945 6883 26979
rect 6825 26939 6883 26945
rect 5169 26911 5227 26917
rect 5169 26877 5181 26911
rect 5215 26908 5227 26911
rect 5258 26908 5264 26920
rect 5215 26880 5264 26908
rect 5215 26877 5227 26880
rect 5169 26871 5227 26877
rect 5258 26868 5264 26880
rect 5316 26868 5322 26920
rect 6730 26868 6736 26920
rect 6788 26908 6794 26920
rect 6840 26908 6868 26939
rect 6914 26936 6920 26988
rect 6972 26936 6978 26988
rect 7190 26936 7196 26988
rect 7248 26936 7254 26988
rect 7377 26979 7435 26985
rect 7377 26945 7389 26979
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 6788 26880 6868 26908
rect 6788 26868 6794 26880
rect 5442 26800 5448 26852
rect 5500 26840 5506 26852
rect 7392 26840 7420 26939
rect 9122 26936 9128 26988
rect 9180 26976 9186 26988
rect 10980 26985 11008 27084
rect 14826 27072 14832 27084
rect 14884 27112 14890 27124
rect 14884 27084 17448 27112
rect 14884 27072 14890 27084
rect 12636 27016 17356 27044
rect 10229 26979 10287 26985
rect 10229 26976 10241 26979
rect 9180 26948 10241 26976
rect 9180 26936 9186 26948
rect 10229 26945 10241 26948
rect 10275 26976 10287 26979
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 10275 26948 10977 26976
rect 10275 26945 10287 26948
rect 10229 26939 10287 26945
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 11974 26936 11980 26988
rect 12032 26976 12038 26988
rect 12636 26985 12664 27016
rect 17328 26985 17356 27016
rect 17420 26985 17448 27084
rect 18966 27004 18972 27056
rect 19024 27004 19030 27056
rect 12621 26979 12679 26985
rect 12621 26976 12633 26979
rect 12032 26948 12633 26976
rect 12032 26936 12038 26948
rect 12621 26945 12633 26948
rect 12667 26945 12679 26979
rect 12621 26939 12679 26945
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 17313 26979 17371 26985
rect 17313 26945 17325 26979
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 12250 26868 12256 26920
rect 12308 26908 12314 26920
rect 13188 26908 13216 26939
rect 12308 26880 13216 26908
rect 17328 26908 17356 26939
rect 17494 26908 17500 26920
rect 17328 26880 17500 26908
rect 12308 26868 12314 26880
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 19702 26868 19708 26920
rect 19760 26868 19766 26920
rect 19978 26868 19984 26920
rect 20036 26868 20042 26920
rect 5500 26812 7420 26840
rect 5500 26800 5506 26812
rect 3602 26732 3608 26784
rect 3660 26772 3666 26784
rect 4433 26775 4491 26781
rect 4433 26772 4445 26775
rect 3660 26744 4445 26772
rect 3660 26732 3666 26744
rect 4433 26741 4445 26744
rect 4479 26741 4491 26775
rect 4433 26735 4491 26741
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26772 7159 26775
rect 7282 26772 7288 26784
rect 7147 26744 7288 26772
rect 7147 26741 7159 26744
rect 7101 26735 7159 26741
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 10318 26732 10324 26784
rect 10376 26732 10382 26784
rect 11057 26775 11115 26781
rect 11057 26741 11069 26775
rect 11103 26772 11115 26775
rect 12066 26772 12072 26784
rect 11103 26744 12072 26772
rect 11103 26741 11115 26744
rect 11057 26735 11115 26741
rect 12066 26732 12072 26744
rect 12124 26732 12130 26784
rect 12710 26732 12716 26784
rect 12768 26732 12774 26784
rect 13078 26732 13084 26784
rect 13136 26732 13142 26784
rect 16206 26732 16212 26784
rect 16264 26772 16270 26784
rect 16669 26775 16727 26781
rect 16669 26772 16681 26775
rect 16264 26744 16681 26772
rect 16264 26732 16270 26744
rect 16669 26741 16681 26744
rect 16715 26741 16727 26775
rect 16669 26735 16727 26741
rect 16850 26732 16856 26784
rect 16908 26772 16914 26784
rect 17497 26775 17555 26781
rect 17497 26772 17509 26775
rect 16908 26744 17509 26772
rect 16908 26732 16914 26744
rect 17497 26741 17509 26744
rect 17543 26741 17555 26775
rect 17497 26735 17555 26741
rect 18138 26732 18144 26784
rect 18196 26772 18202 26784
rect 18233 26775 18291 26781
rect 18233 26772 18245 26775
rect 18196 26744 18245 26772
rect 18196 26732 18202 26744
rect 18233 26741 18245 26744
rect 18279 26741 18291 26775
rect 18233 26735 18291 26741
rect 1104 26682 26864 26704
rect 1104 26630 4169 26682
rect 4221 26630 4233 26682
rect 4285 26630 4297 26682
rect 4349 26630 4361 26682
rect 4413 26630 4425 26682
rect 4477 26630 10608 26682
rect 10660 26630 10672 26682
rect 10724 26630 10736 26682
rect 10788 26630 10800 26682
rect 10852 26630 10864 26682
rect 10916 26630 17047 26682
rect 17099 26630 17111 26682
rect 17163 26630 17175 26682
rect 17227 26630 17239 26682
rect 17291 26630 17303 26682
rect 17355 26630 23486 26682
rect 23538 26630 23550 26682
rect 23602 26630 23614 26682
rect 23666 26630 23678 26682
rect 23730 26630 23742 26682
rect 23794 26630 26864 26682
rect 1104 26608 26864 26630
rect 3786 26528 3792 26580
rect 3844 26568 3850 26580
rect 5442 26568 5448 26580
rect 3844 26540 5448 26568
rect 3844 26528 3850 26540
rect 5442 26528 5448 26540
rect 5500 26528 5506 26580
rect 6825 26571 6883 26577
rect 6825 26537 6837 26571
rect 6871 26568 6883 26571
rect 7190 26568 7196 26580
rect 6871 26540 7196 26568
rect 6871 26537 6883 26540
rect 6825 26531 6883 26537
rect 7190 26528 7196 26540
rect 7248 26528 7254 26580
rect 14366 26528 14372 26580
rect 14424 26577 14430 26580
rect 14424 26571 14473 26577
rect 14424 26537 14427 26571
rect 14461 26568 14473 26571
rect 15979 26571 16037 26577
rect 15979 26568 15991 26571
rect 14461 26540 15991 26568
rect 14461 26537 14473 26540
rect 14424 26531 14473 26537
rect 15979 26537 15991 26540
rect 16025 26537 16037 26571
rect 15979 26531 16037 26537
rect 14424 26528 14430 26531
rect 18966 26528 18972 26580
rect 19024 26528 19030 26580
rect 3605 26503 3663 26509
rect 3605 26469 3617 26503
rect 3651 26500 3663 26503
rect 3651 26472 3832 26500
rect 3651 26469 3663 26472
rect 3605 26463 3663 26469
rect 3804 26432 3832 26472
rect 3878 26460 3884 26512
rect 3936 26500 3942 26512
rect 3936 26472 4108 26500
rect 3936 26460 3942 26472
rect 4080 26441 4108 26472
rect 6472 26472 6684 26500
rect 4065 26435 4123 26441
rect 3804 26404 3924 26432
rect 3326 26324 3332 26376
rect 3384 26324 3390 26376
rect 3602 26324 3608 26376
rect 3660 26324 3666 26376
rect 3786 26324 3792 26376
rect 3844 26324 3850 26376
rect 3896 26296 3924 26404
rect 4065 26401 4077 26435
rect 4111 26432 4123 26435
rect 6472 26432 6500 26472
rect 6656 26444 6684 26472
rect 8110 26460 8116 26512
rect 8168 26500 8174 26512
rect 8665 26503 8723 26509
rect 8665 26500 8677 26503
rect 8168 26472 8677 26500
rect 8168 26460 8174 26472
rect 8665 26469 8677 26472
rect 8711 26469 8723 26503
rect 8665 26463 8723 26469
rect 15838 26460 15844 26512
rect 15896 26460 15902 26512
rect 4111 26404 6500 26432
rect 6549 26435 6607 26441
rect 4111 26401 4123 26404
rect 4065 26395 4123 26401
rect 6549 26401 6561 26435
rect 6595 26401 6607 26435
rect 6549 26395 6607 26401
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 4433 26367 4491 26373
rect 4433 26364 4445 26367
rect 4080 26336 4445 26364
rect 4080 26296 4108 26336
rect 4433 26333 4445 26336
rect 4479 26333 4491 26367
rect 4433 26327 4491 26333
rect 6454 26324 6460 26376
rect 6512 26324 6518 26376
rect 3896 26268 4108 26296
rect 5166 26256 5172 26308
rect 5224 26256 5230 26308
rect 5859 26299 5917 26305
rect 5859 26265 5871 26299
rect 5905 26296 5917 26299
rect 6564 26296 6592 26395
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 6917 26435 6975 26441
rect 6917 26432 6929 26435
rect 6696 26404 6929 26432
rect 6696 26392 6702 26404
rect 6917 26401 6929 26404
rect 6963 26432 6975 26435
rect 6963 26404 11008 26432
rect 6963 26401 6975 26404
rect 6917 26395 6975 26401
rect 10980 26376 11008 26404
rect 13446 26392 13452 26444
rect 13504 26432 13510 26444
rect 15746 26432 15752 26444
rect 13504 26404 13768 26432
rect 13504 26392 13510 26404
rect 7190 26364 7196 26376
rect 7024 26336 7196 26364
rect 7024 26296 7052 26336
rect 7190 26324 7196 26336
rect 7248 26324 7254 26376
rect 7282 26324 7288 26376
rect 7340 26324 7346 26376
rect 9033 26367 9091 26373
rect 9033 26364 9045 26367
rect 8312 26336 9045 26364
rect 5905 26268 6500 26296
rect 6564 26268 7052 26296
rect 8312 26282 8340 26336
rect 9033 26333 9045 26336
rect 9079 26333 9091 26367
rect 9033 26327 9091 26333
rect 9122 26324 9128 26376
rect 9180 26324 9186 26376
rect 10870 26324 10876 26376
rect 10928 26324 10934 26376
rect 10962 26324 10968 26376
rect 11020 26364 11026 26376
rect 11241 26367 11299 26373
rect 11241 26364 11253 26367
rect 11020 26336 11253 26364
rect 11020 26324 11026 26336
rect 11241 26333 11253 26336
rect 11287 26364 11299 26367
rect 11333 26367 11391 26373
rect 11333 26364 11345 26367
rect 11287 26336 11345 26364
rect 11287 26333 11299 26336
rect 11241 26327 11299 26333
rect 11333 26333 11345 26336
rect 11379 26333 11391 26367
rect 11333 26327 11391 26333
rect 12894 26324 12900 26376
rect 12952 26364 12958 26376
rect 13740 26373 13768 26404
rect 13832 26404 15752 26432
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 12952 26336 13553 26364
rect 12952 26324 12958 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26333 13783 26367
rect 13725 26327 13783 26333
rect 9401 26299 9459 26305
rect 5905 26265 5917 26268
rect 5859 26259 5917 26265
rect 3142 26188 3148 26240
rect 3200 26228 3206 26240
rect 3421 26231 3479 26237
rect 3421 26228 3433 26231
rect 3200 26200 3433 26228
rect 3200 26188 3206 26200
rect 3421 26197 3433 26200
rect 3467 26228 3479 26231
rect 3881 26231 3939 26237
rect 3881 26228 3893 26231
rect 3467 26200 3893 26228
rect 3467 26197 3479 26200
rect 3421 26191 3479 26197
rect 3881 26197 3893 26200
rect 3927 26197 3939 26231
rect 6472 26228 6500 26268
rect 9401 26265 9413 26299
rect 9447 26296 9459 26299
rect 9447 26268 9812 26296
rect 9447 26265 9459 26268
rect 9401 26259 9459 26265
rect 7374 26228 7380 26240
rect 6472 26200 7380 26228
rect 3881 26191 3939 26197
rect 7374 26188 7380 26200
rect 7432 26188 7438 26240
rect 9784 26228 9812 26268
rect 10318 26256 10324 26308
rect 10376 26256 10382 26308
rect 11606 26256 11612 26308
rect 11664 26256 11670 26308
rect 12066 26256 12072 26308
rect 12124 26256 12130 26308
rect 13170 26256 13176 26308
rect 13228 26296 13234 26308
rect 13633 26299 13691 26305
rect 13633 26296 13645 26299
rect 13228 26268 13645 26296
rect 13228 26256 13234 26268
rect 13633 26265 13645 26268
rect 13679 26296 13691 26299
rect 13832 26296 13860 26404
rect 15746 26392 15752 26404
rect 15804 26392 15810 26444
rect 16666 26392 16672 26444
rect 16724 26432 16730 26444
rect 17773 26435 17831 26441
rect 17773 26432 17785 26435
rect 16724 26404 17785 26432
rect 16724 26392 16730 26404
rect 17773 26401 17785 26404
rect 17819 26432 17831 26435
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 17819 26404 19257 26432
rect 17819 26401 17831 26404
rect 17773 26395 17831 26401
rect 19245 26401 19257 26404
rect 19291 26432 19303 26435
rect 19978 26432 19984 26444
rect 19291 26404 19984 26432
rect 19291 26401 19303 26404
rect 19245 26395 19303 26401
rect 19978 26392 19984 26404
rect 20036 26392 20042 26444
rect 26142 26392 26148 26444
rect 26200 26392 26206 26444
rect 13909 26367 13967 26373
rect 13909 26333 13921 26367
rect 13955 26333 13967 26367
rect 13909 26327 13967 26333
rect 13679 26268 13860 26296
rect 13924 26296 13952 26327
rect 14090 26324 14096 26376
rect 14148 26324 14154 26376
rect 14274 26324 14280 26376
rect 14332 26324 14338 26376
rect 14458 26324 14464 26376
rect 14516 26364 14522 26376
rect 14553 26367 14611 26373
rect 14553 26364 14565 26367
rect 14516 26336 14565 26364
rect 14516 26324 14522 26336
rect 14553 26333 14565 26336
rect 14599 26333 14611 26367
rect 14553 26327 14611 26333
rect 14826 26324 14832 26376
rect 14884 26324 14890 26376
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26364 15623 26367
rect 16022 26364 16028 26376
rect 15611 26336 16028 26364
rect 15611 26333 15623 26336
rect 15565 26327 15623 26333
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 17402 26324 17408 26376
rect 17460 26324 17466 26376
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26364 18107 26367
rect 18877 26367 18935 26373
rect 18877 26364 18889 26367
rect 18095 26336 18889 26364
rect 18095 26333 18107 26336
rect 18049 26327 18107 26333
rect 18877 26333 18889 26336
rect 18923 26333 18935 26367
rect 18877 26327 18935 26333
rect 15841 26299 15899 26305
rect 15841 26296 15853 26299
rect 13924 26268 15853 26296
rect 13679 26265 13691 26268
rect 13633 26259 13691 26265
rect 15841 26265 15853 26268
rect 15887 26296 15899 26299
rect 16206 26296 16212 26308
rect 15887 26268 16212 26296
rect 15887 26265 15899 26268
rect 15841 26259 15899 26265
rect 16206 26256 16212 26268
rect 16264 26256 16270 26308
rect 16850 26256 16856 26308
rect 16908 26256 16914 26308
rect 18892 26296 18920 26327
rect 25498 26324 25504 26376
rect 25556 26324 25562 26376
rect 18892 26268 19380 26296
rect 19352 26240 19380 26268
rect 19426 26256 19432 26308
rect 19484 26296 19490 26308
rect 19521 26299 19579 26305
rect 19521 26296 19533 26299
rect 19484 26268 19533 26296
rect 19484 26256 19490 26268
rect 19521 26265 19533 26268
rect 19567 26265 19579 26299
rect 19521 26259 19579 26265
rect 19610 26256 19616 26308
rect 19668 26296 19674 26308
rect 19668 26268 20010 26296
rect 19668 26256 19674 26268
rect 21266 26256 21272 26308
rect 21324 26256 21330 26308
rect 10778 26228 10784 26240
rect 9784 26200 10784 26228
rect 10778 26188 10784 26200
rect 10836 26188 10842 26240
rect 12434 26188 12440 26240
rect 12492 26228 12498 26240
rect 13081 26231 13139 26237
rect 13081 26228 13093 26231
rect 12492 26200 13093 26228
rect 12492 26188 12498 26200
rect 13081 26197 13093 26200
rect 13127 26197 13139 26231
rect 13081 26191 13139 26197
rect 13357 26231 13415 26237
rect 13357 26197 13369 26231
rect 13403 26228 13415 26231
rect 13538 26228 13544 26240
rect 13403 26200 13544 26228
rect 13403 26197 13415 26200
rect 13357 26191 13415 26197
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 14093 26231 14151 26237
rect 14093 26228 14105 26231
rect 13872 26200 14105 26228
rect 13872 26188 13878 26200
rect 14093 26197 14105 26200
rect 14139 26197 14151 26231
rect 14093 26191 14151 26197
rect 14734 26188 14740 26240
rect 14792 26188 14798 26240
rect 15657 26231 15715 26237
rect 15657 26197 15669 26231
rect 15703 26228 15715 26231
rect 15746 26228 15752 26240
rect 15703 26200 15752 26228
rect 15703 26197 15715 26200
rect 15657 26191 15715 26197
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 17957 26231 18015 26237
rect 17957 26197 17969 26231
rect 18003 26228 18015 26231
rect 18046 26228 18052 26240
rect 18003 26200 18052 26228
rect 18003 26197 18015 26200
rect 17957 26191 18015 26197
rect 18046 26188 18052 26200
rect 18104 26188 18110 26240
rect 19334 26188 19340 26240
rect 19392 26188 19398 26240
rect 1104 26138 26864 26160
rect 1104 26086 4829 26138
rect 4881 26086 4893 26138
rect 4945 26086 4957 26138
rect 5009 26086 5021 26138
rect 5073 26086 5085 26138
rect 5137 26086 11268 26138
rect 11320 26086 11332 26138
rect 11384 26086 11396 26138
rect 11448 26086 11460 26138
rect 11512 26086 11524 26138
rect 11576 26086 17707 26138
rect 17759 26086 17771 26138
rect 17823 26086 17835 26138
rect 17887 26086 17899 26138
rect 17951 26086 17963 26138
rect 18015 26086 24146 26138
rect 24198 26086 24210 26138
rect 24262 26086 24274 26138
rect 24326 26086 24338 26138
rect 24390 26086 24402 26138
rect 24454 26086 26864 26138
rect 1104 26064 26864 26086
rect 5077 26027 5135 26033
rect 5077 25993 5089 26027
rect 5123 26024 5135 26027
rect 5166 26024 5172 26036
rect 5123 25996 5172 26024
rect 5123 25993 5135 25996
rect 5077 25987 5135 25993
rect 5166 25984 5172 25996
rect 5224 25984 5230 26036
rect 7190 25984 7196 26036
rect 7248 26024 7254 26036
rect 7285 26027 7343 26033
rect 7285 26024 7297 26027
rect 7248 25996 7297 26024
rect 7248 25984 7254 25996
rect 7285 25993 7297 25996
rect 7331 25993 7343 26027
rect 7285 25987 7343 25993
rect 11333 26027 11391 26033
rect 11333 25993 11345 26027
rect 11379 26024 11391 26027
rect 11606 26024 11612 26036
rect 11379 25996 11612 26024
rect 11379 25993 11391 25996
rect 11333 25987 11391 25993
rect 11606 25984 11612 25996
rect 11664 25984 11670 26036
rect 11698 25984 11704 26036
rect 11756 26024 11762 26036
rect 12250 26024 12256 26036
rect 11756 25996 12256 26024
rect 11756 25984 11762 25996
rect 12250 25984 12256 25996
rect 12308 25984 12314 26036
rect 13814 26024 13820 26036
rect 13280 25996 13820 26024
rect 4801 25959 4859 25965
rect 4801 25956 4813 25959
rect 4186 25928 4813 25956
rect 4801 25925 4813 25928
rect 4847 25925 4859 25959
rect 4801 25919 4859 25925
rect 6454 25916 6460 25968
rect 6512 25956 6518 25968
rect 7098 25956 7104 25968
rect 6512 25928 7104 25956
rect 6512 25916 6518 25928
rect 7098 25916 7104 25928
rect 7156 25916 7162 25968
rect 7374 25916 7380 25968
rect 7432 25956 7438 25968
rect 7432 25928 7972 25956
rect 7432 25916 7438 25928
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25857 2835 25891
rect 2777 25851 2835 25857
rect 2792 25820 2820 25851
rect 3142 25848 3148 25900
rect 3200 25848 3206 25900
rect 4893 25891 4951 25897
rect 4893 25857 4905 25891
rect 4939 25888 4951 25891
rect 4985 25891 5043 25897
rect 4985 25888 4997 25891
rect 4939 25860 4997 25888
rect 4939 25857 4951 25860
rect 4893 25851 4951 25857
rect 4985 25857 4997 25860
rect 5031 25888 5043 25891
rect 5994 25888 6000 25900
rect 5031 25860 6000 25888
rect 5031 25857 5043 25860
rect 4985 25851 5043 25857
rect 5994 25848 6000 25860
rect 6052 25848 6058 25900
rect 7009 25891 7067 25897
rect 7009 25857 7021 25891
rect 7055 25888 7067 25891
rect 7116 25888 7144 25916
rect 7055 25860 7144 25888
rect 7469 25891 7527 25897
rect 7055 25857 7067 25860
rect 7009 25851 7067 25857
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7558 25888 7564 25900
rect 7515 25860 7564 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7558 25848 7564 25860
rect 7616 25888 7622 25900
rect 7944 25897 7972 25928
rect 9674 25916 9680 25968
rect 9732 25916 9738 25968
rect 10962 25956 10968 25968
rect 10428 25928 10968 25956
rect 10428 25897 10456 25928
rect 10962 25916 10968 25928
rect 11020 25916 11026 25968
rect 11974 25956 11980 25968
rect 11072 25928 11980 25956
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 7616 25860 7757 25888
rect 7616 25848 7622 25860
rect 7745 25857 7757 25860
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 2958 25820 2964 25832
rect 2792 25792 2964 25820
rect 2958 25780 2964 25792
rect 3016 25820 3022 25832
rect 3878 25820 3884 25832
rect 3016 25792 3884 25820
rect 3016 25780 3022 25792
rect 3878 25780 3884 25792
rect 3936 25780 3942 25832
rect 7101 25823 7159 25829
rect 7101 25789 7113 25823
rect 7147 25789 7159 25823
rect 7101 25783 7159 25789
rect 7006 25712 7012 25764
rect 7064 25752 7070 25764
rect 7116 25752 7144 25783
rect 7374 25780 7380 25832
rect 7432 25820 7438 25832
rect 7653 25823 7711 25829
rect 7653 25820 7665 25823
rect 7432 25792 7665 25820
rect 7432 25780 7438 25792
rect 7653 25789 7665 25792
rect 7699 25789 7711 25823
rect 7760 25820 7788 25851
rect 10778 25848 10784 25900
rect 10836 25888 10842 25900
rect 11072 25897 11100 25928
rect 11974 25916 11980 25928
rect 12032 25916 12038 25968
rect 12158 25965 12164 25968
rect 12115 25959 12164 25965
rect 12115 25925 12127 25959
rect 12161 25925 12164 25959
rect 12115 25919 12164 25925
rect 12158 25916 12164 25919
rect 12216 25916 12222 25968
rect 11057 25891 11115 25897
rect 10836 25860 11008 25888
rect 10836 25848 10842 25860
rect 10980 25832 11008 25860
rect 11057 25857 11069 25891
rect 11103 25857 11115 25891
rect 11057 25851 11115 25857
rect 11790 25848 11796 25900
rect 11848 25848 11854 25900
rect 11885 25891 11943 25897
rect 11885 25857 11897 25891
rect 11931 25857 11943 25891
rect 12253 25891 12311 25897
rect 12253 25878 12265 25891
rect 11885 25851 11943 25857
rect 12130 25857 12265 25878
rect 12299 25857 12311 25891
rect 12130 25851 12311 25857
rect 8619 25823 8677 25829
rect 8619 25820 8631 25823
rect 7760 25792 8631 25820
rect 7653 25783 7711 25789
rect 8619 25789 8631 25792
rect 8665 25789 8677 25823
rect 8619 25783 8677 25789
rect 10045 25823 10103 25829
rect 10045 25789 10057 25823
rect 10091 25820 10103 25823
rect 10226 25820 10232 25832
rect 10091 25792 10232 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10226 25780 10232 25792
rect 10284 25780 10290 25832
rect 10873 25823 10931 25829
rect 10873 25789 10885 25823
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 7745 25755 7803 25761
rect 7745 25752 7757 25755
rect 7064 25724 7757 25752
rect 7064 25712 7070 25724
rect 7745 25721 7757 25724
rect 7791 25721 7803 25755
rect 10888 25752 10916 25783
rect 10962 25780 10968 25832
rect 11020 25780 11026 25832
rect 11149 25823 11207 25829
rect 11149 25789 11161 25823
rect 11195 25820 11207 25823
rect 11698 25820 11704 25832
rect 11195 25792 11704 25820
rect 11195 25789 11207 25792
rect 11149 25783 11207 25789
rect 11698 25780 11704 25792
rect 11756 25780 11762 25832
rect 11900 25820 11928 25851
rect 12130 25850 12296 25851
rect 12130 25832 12158 25850
rect 12342 25848 12348 25900
rect 12400 25848 12406 25900
rect 12434 25848 12440 25900
rect 12492 25848 12498 25900
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 13280 25888 13308 25996
rect 13814 25984 13820 25996
rect 13872 25984 13878 26036
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 18463 26027 18521 26033
rect 18463 26024 18475 26027
rect 17552 25996 18475 26024
rect 17552 25984 17558 25996
rect 18463 25993 18475 25996
rect 18509 25993 18521 26027
rect 18463 25987 18521 25993
rect 19610 25984 19616 26036
rect 19668 25984 19674 26036
rect 14734 25916 14740 25968
rect 14792 25916 14798 25968
rect 15838 25916 15844 25968
rect 15896 25956 15902 25968
rect 16301 25959 16359 25965
rect 16301 25956 16313 25959
rect 15896 25928 16313 25956
rect 15896 25916 15902 25928
rect 16301 25925 16313 25928
rect 16347 25925 16359 25959
rect 16301 25919 16359 25925
rect 18046 25916 18052 25968
rect 18104 25916 18110 25968
rect 12575 25860 13308 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 15746 25848 15752 25900
rect 15804 25848 15810 25900
rect 15930 25848 15936 25900
rect 15988 25848 15994 25900
rect 16022 25848 16028 25900
rect 16080 25848 16086 25900
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16163 25860 17049 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 11974 25820 11980 25832
rect 11900 25792 11980 25820
rect 11974 25780 11980 25792
rect 12032 25780 12038 25832
rect 12066 25780 12072 25832
rect 12124 25792 12158 25832
rect 12452 25820 12480 25848
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 12452 25792 12633 25820
rect 12124 25780 12130 25792
rect 12621 25789 12633 25792
rect 12667 25789 12679 25823
rect 12621 25783 12679 25789
rect 13354 25780 13360 25832
rect 13412 25780 13418 25832
rect 13538 25780 13544 25832
rect 13596 25820 13602 25832
rect 13725 25823 13783 25829
rect 13725 25820 13737 25823
rect 13596 25792 13737 25820
rect 13596 25780 13602 25792
rect 13725 25789 13737 25792
rect 13771 25789 13783 25823
rect 13725 25783 13783 25789
rect 11514 25752 11520 25764
rect 10888 25724 11520 25752
rect 7745 25715 7803 25721
rect 11514 25712 11520 25724
rect 11572 25712 11578 25764
rect 12437 25755 12495 25761
rect 12437 25721 12449 25755
rect 12483 25752 12495 25755
rect 12894 25752 12900 25764
rect 12483 25724 12900 25752
rect 12483 25721 12495 25724
rect 12437 25715 12495 25721
rect 12894 25712 12900 25724
rect 12952 25712 12958 25764
rect 15933 25755 15991 25761
rect 15933 25721 15945 25755
rect 15979 25752 15991 25755
rect 16316 25752 16344 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19392 25860 19533 25888
rect 19392 25848 19398 25860
rect 19521 25857 19533 25860
rect 19567 25888 19579 25891
rect 20162 25888 20168 25900
rect 19567 25860 20168 25888
rect 19567 25857 19579 25860
rect 19521 25851 19579 25857
rect 20162 25848 20168 25860
rect 20220 25848 20226 25900
rect 16666 25780 16672 25832
rect 16724 25780 16730 25832
rect 15979 25724 16344 25752
rect 15979 25721 15991 25724
rect 15933 25715 15991 25721
rect 4571 25687 4629 25693
rect 4571 25653 4583 25687
rect 4617 25684 4629 25687
rect 5258 25684 5264 25696
rect 4617 25656 5264 25684
rect 4617 25653 4629 25656
rect 4571 25647 4629 25653
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 6641 25687 6699 25693
rect 6641 25653 6653 25687
rect 6687 25684 6699 25687
rect 6914 25684 6920 25696
rect 6687 25656 6920 25684
rect 6687 25653 6699 25656
rect 6641 25647 6699 25653
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 11054 25644 11060 25696
rect 11112 25684 11118 25696
rect 11609 25687 11667 25693
rect 11609 25684 11621 25687
rect 11112 25656 11621 25684
rect 11112 25644 11118 25656
rect 11609 25653 11621 25656
rect 11655 25653 11667 25687
rect 11609 25647 11667 25653
rect 12986 25644 12992 25696
rect 13044 25684 13050 25696
rect 13265 25687 13323 25693
rect 13265 25684 13277 25687
rect 13044 25656 13277 25684
rect 13044 25644 13050 25656
rect 13265 25653 13277 25656
rect 13311 25653 13323 25687
rect 13265 25647 13323 25653
rect 14090 25644 14096 25696
rect 14148 25684 14154 25696
rect 14550 25684 14556 25696
rect 14148 25656 14556 25684
rect 14148 25644 14154 25656
rect 14550 25644 14556 25656
rect 14608 25684 14614 25696
rect 15151 25687 15209 25693
rect 15151 25684 15163 25687
rect 14608 25656 15163 25684
rect 14608 25644 14614 25656
rect 15151 25653 15163 25656
rect 15197 25653 15209 25687
rect 15151 25647 15209 25653
rect 16301 25687 16359 25693
rect 16301 25653 16313 25687
rect 16347 25684 16359 25687
rect 17402 25684 17408 25696
rect 16347 25656 17408 25684
rect 16347 25653 16359 25656
rect 16301 25647 16359 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 1104 25594 26864 25616
rect 1104 25542 4169 25594
rect 4221 25542 4233 25594
rect 4285 25542 4297 25594
rect 4349 25542 4361 25594
rect 4413 25542 4425 25594
rect 4477 25542 10608 25594
rect 10660 25542 10672 25594
rect 10724 25542 10736 25594
rect 10788 25542 10800 25594
rect 10852 25542 10864 25594
rect 10916 25542 17047 25594
rect 17099 25542 17111 25594
rect 17163 25542 17175 25594
rect 17227 25542 17239 25594
rect 17291 25542 17303 25594
rect 17355 25542 23486 25594
rect 23538 25542 23550 25594
rect 23602 25542 23614 25594
rect 23666 25542 23678 25594
rect 23730 25542 23742 25594
rect 23794 25542 26864 25594
rect 1104 25520 26864 25542
rect 4522 25440 4528 25492
rect 4580 25480 4586 25492
rect 4617 25483 4675 25489
rect 4617 25480 4629 25483
rect 4580 25452 4629 25480
rect 4580 25440 4586 25452
rect 4617 25449 4629 25452
rect 4663 25449 4675 25483
rect 4617 25443 4675 25449
rect 7098 25440 7104 25492
rect 7156 25440 7162 25492
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 9732 25452 9965 25480
rect 9732 25440 9738 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 9953 25443 10011 25449
rect 11514 25440 11520 25492
rect 11572 25440 11578 25492
rect 12066 25480 12072 25492
rect 11716 25452 12072 25480
rect 4433 25415 4491 25421
rect 4433 25381 4445 25415
rect 4479 25412 4491 25415
rect 5442 25412 5448 25424
rect 4479 25384 5448 25412
rect 4479 25381 4491 25384
rect 4433 25375 4491 25381
rect 5442 25372 5448 25384
rect 5500 25372 5506 25424
rect 5994 25372 6000 25424
rect 6052 25412 6058 25424
rect 9122 25412 9128 25424
rect 6052 25384 9128 25412
rect 6052 25372 6058 25384
rect 9122 25372 9128 25384
rect 9180 25372 9186 25424
rect 11425 25415 11483 25421
rect 11425 25381 11437 25415
rect 11471 25412 11483 25415
rect 11716 25412 11744 25452
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12158 25440 12164 25492
rect 12216 25480 12222 25492
rect 12253 25483 12311 25489
rect 12253 25480 12265 25483
rect 12216 25452 12265 25480
rect 12216 25440 12222 25452
rect 12253 25449 12265 25452
rect 12299 25480 12311 25483
rect 13170 25480 13176 25492
rect 12299 25452 13176 25480
rect 12299 25449 12311 25452
rect 12253 25443 12311 25449
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 13354 25440 13360 25492
rect 13412 25480 13418 25492
rect 13412 25452 13860 25480
rect 13412 25440 13418 25452
rect 12342 25412 12348 25424
rect 11471 25384 11744 25412
rect 11900 25384 12348 25412
rect 11471 25381 11483 25384
rect 11425 25375 11483 25381
rect 4062 25304 4068 25356
rect 4120 25304 4126 25356
rect 9140 25344 9168 25372
rect 11900 25353 11928 25384
rect 12342 25372 12348 25384
rect 12400 25412 12406 25424
rect 12621 25415 12679 25421
rect 12621 25412 12633 25415
rect 12400 25384 12633 25412
rect 12400 25372 12406 25384
rect 12621 25381 12633 25384
rect 12667 25412 12679 25415
rect 13449 25415 13507 25421
rect 13449 25412 13461 25415
rect 12667 25384 13461 25412
rect 12667 25381 12679 25384
rect 12621 25375 12679 25381
rect 13449 25381 13461 25384
rect 13495 25381 13507 25415
rect 13832 25412 13860 25452
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 14458 25480 14464 25492
rect 13964 25452 14464 25480
rect 13964 25440 13970 25452
rect 14458 25440 14464 25452
rect 14516 25440 14522 25492
rect 15473 25483 15531 25489
rect 15473 25449 15485 25483
rect 15519 25480 15531 25483
rect 16022 25480 16028 25492
rect 15519 25452 16028 25480
rect 15519 25449 15531 25452
rect 15473 25443 15531 25449
rect 16022 25440 16028 25452
rect 16080 25440 16086 25492
rect 19702 25440 19708 25492
rect 19760 25480 19766 25492
rect 19797 25483 19855 25489
rect 19797 25480 19809 25483
rect 19760 25452 19809 25480
rect 19760 25440 19766 25452
rect 19797 25449 19809 25452
rect 19843 25449 19855 25483
rect 19797 25443 19855 25449
rect 16666 25412 16672 25424
rect 13832 25384 16672 25412
rect 13449 25375 13507 25381
rect 16666 25372 16672 25384
rect 16724 25412 16730 25424
rect 16942 25412 16948 25424
rect 16724 25384 16948 25412
rect 16724 25372 16730 25384
rect 16942 25372 16948 25384
rect 17000 25372 17006 25424
rect 18506 25372 18512 25424
rect 18564 25412 18570 25424
rect 18564 25384 18644 25412
rect 18564 25372 18570 25384
rect 9769 25347 9827 25353
rect 9140 25316 9260 25344
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25276 4031 25279
rect 4522 25276 4528 25288
rect 4019 25248 4528 25276
rect 4019 25245 4031 25248
rect 3973 25239 4031 25245
rect 4522 25236 4528 25248
rect 4580 25236 4586 25288
rect 4893 25279 4951 25285
rect 4893 25245 4905 25279
rect 4939 25276 4951 25279
rect 5258 25276 5264 25288
rect 4939 25248 5264 25276
rect 4939 25245 4951 25248
rect 4893 25239 4951 25245
rect 5258 25236 5264 25248
rect 5316 25236 5322 25288
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25276 6883 25279
rect 6871 25248 6905 25276
rect 6871 25245 6883 25248
rect 6825 25239 6883 25245
rect 3602 25168 3608 25220
rect 3660 25208 3666 25220
rect 4706 25208 4712 25220
rect 3660 25180 4712 25208
rect 3660 25168 3666 25180
rect 4706 25168 4712 25180
rect 4764 25208 4770 25220
rect 4801 25211 4859 25217
rect 4801 25208 4813 25211
rect 4764 25180 4813 25208
rect 4764 25168 4770 25180
rect 4801 25177 4813 25180
rect 4847 25177 4859 25211
rect 6840 25208 6868 25239
rect 7650 25236 7656 25288
rect 7708 25276 7714 25288
rect 9125 25279 9183 25285
rect 9125 25276 9137 25279
rect 7708 25248 9137 25276
rect 7708 25236 7714 25248
rect 9125 25245 9137 25248
rect 9171 25245 9183 25279
rect 9232 25276 9260 25316
rect 9769 25313 9781 25347
rect 9815 25344 9827 25347
rect 11149 25347 11207 25353
rect 9815 25316 10180 25344
rect 9815 25313 9827 25316
rect 9769 25307 9827 25313
rect 10152 25285 10180 25316
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 11885 25347 11943 25353
rect 11885 25344 11897 25347
rect 11195 25316 11897 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 11885 25313 11897 25316
rect 11931 25313 11943 25347
rect 11885 25307 11943 25313
rect 13722 25304 13728 25356
rect 13780 25344 13786 25356
rect 13817 25347 13875 25353
rect 13817 25344 13829 25347
rect 13780 25316 13829 25344
rect 13780 25304 13786 25316
rect 13817 25313 13829 25316
rect 13863 25344 13875 25347
rect 14366 25344 14372 25356
rect 13863 25316 14372 25344
rect 13863 25313 13875 25316
rect 13817 25307 13875 25313
rect 14366 25304 14372 25316
rect 14424 25344 14430 25356
rect 18616 25353 18644 25384
rect 14921 25347 14979 25353
rect 14424 25316 14872 25344
rect 14424 25304 14430 25316
rect 10045 25279 10103 25285
rect 10045 25276 10057 25279
rect 9232 25248 10057 25276
rect 9125 25239 9183 25245
rect 10045 25245 10057 25248
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 10962 25236 10968 25288
rect 11020 25276 11026 25288
rect 11057 25279 11115 25285
rect 11057 25276 11069 25279
rect 11020 25248 11069 25276
rect 11020 25236 11026 25248
rect 11057 25245 11069 25248
rect 11103 25276 11115 25279
rect 11103 25270 11652 25276
rect 11698 25270 11704 25288
rect 11103 25248 11704 25270
rect 11103 25245 11115 25248
rect 11057 25239 11115 25245
rect 11624 25242 11704 25248
rect 11698 25236 11704 25242
rect 11756 25236 11762 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25245 11851 25279
rect 11793 25239 11851 25245
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25245 12035 25279
rect 11977 25239 12035 25245
rect 7085 25211 7143 25217
rect 4801 25171 4859 25177
rect 4908 25180 6960 25208
rect 4338 25100 4344 25152
rect 4396 25100 4402 25152
rect 4614 25149 4620 25152
rect 4601 25143 4620 25149
rect 4601 25109 4613 25143
rect 4672 25140 4678 25152
rect 4908 25140 4936 25180
rect 4672 25112 4936 25140
rect 4985 25143 5043 25149
rect 4601 25103 4620 25109
rect 4614 25100 4620 25103
rect 4672 25100 4678 25112
rect 4985 25109 4997 25143
rect 5031 25140 5043 25143
rect 5166 25140 5172 25152
rect 5031 25112 5172 25140
rect 5031 25109 5043 25112
rect 4985 25103 5043 25109
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 6733 25143 6791 25149
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 6822 25140 6828 25152
rect 6779 25112 6828 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 6932 25149 6960 25180
rect 7085 25177 7097 25211
rect 7131 25208 7143 25211
rect 7190 25208 7196 25220
rect 7131 25180 7196 25208
rect 7131 25177 7143 25180
rect 7085 25171 7143 25177
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 7285 25211 7343 25217
rect 7285 25177 7297 25211
rect 7331 25208 7343 25211
rect 7374 25208 7380 25220
rect 7331 25180 7380 25208
rect 7331 25177 7343 25180
rect 7285 25171 7343 25177
rect 7374 25168 7380 25180
rect 7432 25168 7438 25220
rect 11808 25208 11836 25239
rect 11882 25208 11888 25220
rect 11808 25180 11888 25208
rect 11882 25168 11888 25180
rect 11940 25168 11946 25220
rect 6917 25143 6975 25149
rect 6917 25109 6929 25143
rect 6963 25109 6975 25143
rect 6917 25103 6975 25109
rect 10226 25100 10232 25152
rect 10284 25100 10290 25152
rect 11992 25140 12020 25239
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 12710 25236 12716 25288
rect 12768 25236 12774 25288
rect 13538 25236 13544 25288
rect 13596 25276 13602 25288
rect 13633 25279 13691 25285
rect 13633 25276 13645 25279
rect 13596 25248 13645 25276
rect 13596 25236 13602 25248
rect 13633 25245 13645 25248
rect 13679 25245 13691 25279
rect 13633 25239 13691 25245
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14550 25236 14556 25288
rect 14608 25236 14614 25288
rect 14844 25285 14872 25316
rect 14921 25313 14933 25347
rect 14967 25344 14979 25347
rect 15657 25347 15715 25353
rect 14967 25316 15332 25344
rect 14967 25313 14979 25316
rect 14921 25307 14979 25313
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25276 15071 25279
rect 15194 25276 15200 25288
rect 15059 25248 15200 25276
rect 15059 25245 15071 25248
rect 15013 25239 15071 25245
rect 13909 25211 13967 25217
rect 13909 25177 13921 25211
rect 13955 25208 13967 25211
rect 14292 25208 14320 25236
rect 15028 25208 15056 25239
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 15304 25285 15332 25316
rect 15657 25313 15669 25347
rect 15703 25313 15715 25347
rect 15657 25307 15715 25313
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 18601 25347 18659 25353
rect 16163 25316 16620 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25276 15347 25279
rect 15672 25276 15700 25307
rect 15335 25248 15700 25276
rect 15749 25279 15807 25285
rect 15335 25245 15347 25248
rect 15289 25239 15347 25245
rect 15749 25245 15761 25279
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 13955 25180 15056 25208
rect 13955 25177 13967 25180
rect 13909 25171 13967 25177
rect 15102 25168 15108 25220
rect 15160 25168 15166 25220
rect 15654 25168 15660 25220
rect 15712 25208 15718 25220
rect 15764 25208 15792 25239
rect 16206 25236 16212 25288
rect 16264 25236 16270 25288
rect 16592 25285 16620 25316
rect 18601 25313 18613 25347
rect 18647 25313 18659 25347
rect 18601 25307 18659 25313
rect 16577 25279 16635 25285
rect 16577 25245 16589 25279
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18555 25248 18644 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18616 25220 18644 25248
rect 19334 25236 19340 25288
rect 19392 25236 19398 25288
rect 19429 25279 19487 25285
rect 19429 25245 19441 25279
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 15712 25180 15792 25208
rect 15712 25168 15718 25180
rect 16390 25168 16396 25220
rect 16448 25168 16454 25220
rect 16485 25211 16543 25217
rect 16485 25177 16497 25211
rect 16531 25177 16543 25211
rect 16485 25171 16543 25177
rect 12434 25140 12440 25152
rect 11992 25112 12440 25140
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 14090 25100 14096 25152
rect 14148 25100 14154 25152
rect 15746 25100 15752 25152
rect 15804 25140 15810 25152
rect 16500 25140 16528 25171
rect 18598 25168 18604 25220
rect 18656 25208 18662 25220
rect 19444 25208 19472 25239
rect 19518 25236 19524 25288
rect 19576 25236 19582 25288
rect 19610 25236 19616 25288
rect 19668 25236 19674 25288
rect 18656 25180 19472 25208
rect 18656 25168 18662 25180
rect 15804 25112 16528 25140
rect 16761 25143 16819 25149
rect 15804 25100 15810 25112
rect 16761 25109 16773 25143
rect 16807 25140 16819 25143
rect 16850 25140 16856 25152
rect 16807 25112 16856 25140
rect 16807 25109 16819 25112
rect 16761 25103 16819 25109
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 18782 25100 18788 25152
rect 18840 25140 18846 25152
rect 18877 25143 18935 25149
rect 18877 25140 18889 25143
rect 18840 25112 18889 25140
rect 18840 25100 18846 25112
rect 18877 25109 18889 25112
rect 18923 25109 18935 25143
rect 18877 25103 18935 25109
rect 1104 25050 26864 25072
rect 1104 24998 4829 25050
rect 4881 24998 4893 25050
rect 4945 24998 4957 25050
rect 5009 24998 5021 25050
rect 5073 24998 5085 25050
rect 5137 24998 11268 25050
rect 11320 24998 11332 25050
rect 11384 24998 11396 25050
rect 11448 24998 11460 25050
rect 11512 24998 11524 25050
rect 11576 24998 17707 25050
rect 17759 24998 17771 25050
rect 17823 24998 17835 25050
rect 17887 24998 17899 25050
rect 17951 24998 17963 25050
rect 18015 24998 24146 25050
rect 24198 24998 24210 25050
rect 24262 24998 24274 25050
rect 24326 24998 24338 25050
rect 24390 24998 24402 25050
rect 24454 24998 26864 25050
rect 1104 24976 26864 24998
rect 4430 24896 4436 24948
rect 4488 24936 4494 24948
rect 4525 24939 4583 24945
rect 4525 24936 4537 24939
rect 4488 24908 4537 24936
rect 4488 24896 4494 24908
rect 4525 24905 4537 24908
rect 4571 24936 4583 24939
rect 6730 24936 6736 24948
rect 4571 24908 6736 24936
rect 4571 24905 4583 24908
rect 4525 24899 4583 24905
rect 6730 24896 6736 24908
rect 6788 24896 6794 24948
rect 11790 24896 11796 24948
rect 11848 24936 11854 24948
rect 11885 24939 11943 24945
rect 11885 24936 11897 24939
rect 11848 24908 11897 24936
rect 11848 24896 11854 24908
rect 11885 24905 11897 24908
rect 11931 24905 11943 24939
rect 11885 24899 11943 24905
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 12345 24939 12403 24945
rect 12345 24936 12357 24939
rect 12032 24908 12357 24936
rect 12032 24896 12038 24908
rect 12345 24905 12357 24908
rect 12391 24905 12403 24939
rect 12345 24899 12403 24905
rect 12802 24896 12808 24948
rect 12860 24936 12866 24948
rect 13538 24936 13544 24948
rect 12860 24908 13544 24936
rect 12860 24896 12866 24908
rect 13538 24896 13544 24908
rect 13596 24936 13602 24948
rect 14550 24936 14556 24948
rect 13596 24908 14556 24936
rect 13596 24896 13602 24908
rect 3142 24828 3148 24880
rect 3200 24828 3206 24880
rect 4249 24871 4307 24877
rect 4249 24837 4261 24871
rect 4295 24868 4307 24871
rect 4338 24868 4344 24880
rect 4295 24840 4344 24868
rect 4295 24837 4307 24840
rect 4249 24831 4307 24837
rect 4338 24828 4344 24840
rect 4396 24828 4402 24880
rect 4614 24828 4620 24880
rect 4672 24868 4678 24880
rect 5074 24868 5080 24880
rect 4672 24840 5080 24868
rect 4672 24828 4678 24840
rect 5074 24828 5080 24840
rect 5132 24828 5138 24880
rect 6748 24868 6776 24896
rect 6656 24840 6776 24868
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 1765 24803 1823 24809
rect 1765 24800 1777 24803
rect 1452 24772 1777 24800
rect 1452 24760 1458 24772
rect 1765 24769 1777 24772
rect 1811 24800 1823 24803
rect 1811 24772 2268 24800
rect 1811 24769 1823 24772
rect 1765 24763 1823 24769
rect 2133 24735 2191 24741
rect 2133 24732 2145 24735
rect 1780 24704 2145 24732
rect 1780 24596 1808 24704
rect 2133 24701 2145 24704
rect 2179 24701 2191 24735
rect 2240 24732 2268 24772
rect 3970 24760 3976 24812
rect 4028 24760 4034 24812
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4120 24772 4476 24800
rect 4120 24760 4126 24772
rect 2958 24732 2964 24744
rect 2240 24704 2964 24732
rect 2133 24695 2191 24701
rect 2958 24692 2964 24704
rect 3016 24692 3022 24744
rect 3878 24692 3884 24744
rect 3936 24692 3942 24744
rect 4338 24692 4344 24744
rect 4396 24692 4402 24744
rect 4448 24732 4476 24772
rect 4706 24760 4712 24812
rect 4764 24760 4770 24812
rect 4798 24760 4804 24812
rect 4856 24760 4862 24812
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24800 5043 24803
rect 5166 24800 5172 24812
rect 5031 24772 5172 24800
rect 5031 24769 5043 24772
rect 4985 24763 5043 24769
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 5258 24760 5264 24812
rect 5316 24800 5322 24812
rect 5445 24803 5503 24809
rect 5445 24800 5457 24803
rect 5316 24772 5457 24800
rect 5316 24760 5322 24772
rect 5445 24769 5457 24772
rect 5491 24769 5503 24803
rect 5445 24763 5503 24769
rect 5997 24803 6055 24809
rect 5997 24769 6009 24803
rect 6043 24769 6055 24803
rect 5997 24763 6055 24769
rect 4448 24704 4936 24732
rect 4908 24673 4936 24704
rect 5074 24692 5080 24744
rect 5132 24732 5138 24744
rect 5353 24735 5411 24741
rect 5353 24732 5365 24735
rect 5132 24704 5365 24732
rect 5132 24692 5138 24704
rect 5353 24701 5365 24704
rect 5399 24701 5411 24735
rect 5353 24695 5411 24701
rect 5534 24692 5540 24744
rect 5592 24692 5598 24744
rect 5626 24692 5632 24744
rect 5684 24692 5690 24744
rect 4893 24667 4951 24673
rect 3436 24636 4660 24664
rect 3436 24596 3464 24636
rect 3602 24605 3608 24608
rect 1780 24568 3464 24596
rect 3559 24599 3608 24605
rect 3559 24565 3571 24599
rect 3605 24565 3608 24599
rect 3559 24559 3608 24565
rect 3602 24556 3608 24559
rect 3660 24556 3666 24608
rect 3694 24556 3700 24608
rect 3752 24556 3758 24608
rect 4632 24596 4660 24636
rect 4893 24633 4905 24667
rect 4939 24664 4951 24667
rect 6012 24664 6040 24763
rect 6178 24760 6184 24812
rect 6236 24760 6242 24812
rect 6362 24760 6368 24812
rect 6420 24760 6426 24812
rect 6546 24760 6552 24812
rect 6604 24760 6610 24812
rect 6656 24809 6684 24840
rect 11698 24828 11704 24880
rect 11756 24868 11762 24880
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 11756 24840 12081 24868
rect 11756 24828 11762 24840
rect 12069 24837 12081 24840
rect 12115 24868 12127 24871
rect 13709 24871 13767 24877
rect 12115 24840 12434 24868
rect 12115 24837 12127 24840
rect 12069 24831 12127 24837
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24769 6699 24803
rect 6641 24763 6699 24769
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24769 6791 24803
rect 6733 24763 6791 24769
rect 6089 24735 6147 24741
rect 6089 24701 6101 24735
rect 6135 24732 6147 24735
rect 6748 24732 6776 24763
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 7650 24760 7656 24812
rect 7708 24800 7714 24812
rect 7929 24803 7987 24809
rect 7929 24800 7941 24803
rect 7708 24772 7941 24800
rect 7708 24760 7714 24772
rect 7929 24769 7941 24772
rect 7975 24769 7987 24803
rect 7929 24763 7987 24769
rect 12250 24760 12256 24812
rect 12308 24760 12314 24812
rect 6135 24704 6776 24732
rect 6135 24701 6147 24704
rect 6089 24695 6147 24701
rect 7006 24692 7012 24744
rect 7064 24732 7070 24744
rect 7484 24732 7512 24760
rect 8018 24732 8024 24744
rect 7064 24704 8024 24732
rect 7064 24692 7070 24704
rect 8018 24692 8024 24704
rect 8076 24692 8082 24744
rect 8110 24692 8116 24744
rect 8168 24692 8174 24744
rect 8202 24692 8208 24744
rect 8260 24692 8266 24744
rect 12406 24732 12434 24840
rect 12820 24840 13124 24868
rect 12621 24803 12679 24809
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 12820 24800 12848 24840
rect 13096 24812 13124 24840
rect 13709 24837 13721 24871
rect 13755 24868 13767 24871
rect 13814 24868 13820 24880
rect 13755 24840 13820 24868
rect 13755 24837 13767 24840
rect 13709 24831 13767 24837
rect 13814 24828 13820 24840
rect 13872 24828 13878 24880
rect 13924 24877 13952 24908
rect 14550 24896 14556 24908
rect 14608 24896 14614 24948
rect 16117 24939 16175 24945
rect 16117 24905 16129 24939
rect 16163 24936 16175 24939
rect 16390 24936 16396 24948
rect 16163 24908 16396 24936
rect 16163 24905 16175 24908
rect 16117 24899 16175 24905
rect 16390 24896 16396 24908
rect 16448 24896 16454 24948
rect 13909 24871 13967 24877
rect 13909 24837 13921 24871
rect 13955 24837 13967 24871
rect 13909 24831 13967 24837
rect 14458 24828 14464 24880
rect 14516 24868 14522 24880
rect 15654 24868 15660 24880
rect 14516 24840 15660 24868
rect 14516 24828 14522 24840
rect 12667 24772 12848 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 12894 24760 12900 24812
rect 12952 24760 12958 24812
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 12526 24732 12532 24744
rect 12406 24704 12532 24732
rect 12526 24692 12532 24704
rect 12584 24732 12590 24744
rect 12912 24732 12940 24760
rect 12584 24704 12940 24732
rect 13004 24732 13032 24763
rect 13078 24760 13084 24812
rect 13136 24760 13142 24812
rect 13262 24760 13268 24812
rect 13320 24760 13326 24812
rect 13446 24760 13452 24812
rect 13504 24760 13510 24812
rect 13832 24800 13860 24828
rect 15212 24809 15240 24840
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 15930 24828 15936 24880
rect 15988 24828 15994 24880
rect 19352 24840 19564 24868
rect 15197 24803 15255 24809
rect 13832 24772 14504 24800
rect 14090 24732 14096 24744
rect 13004 24704 14096 24732
rect 12584 24692 12590 24704
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 14476 24732 14504 24772
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15749 24803 15807 24809
rect 15749 24800 15761 24803
rect 15197 24763 15255 24769
rect 15580 24772 15761 24800
rect 15102 24732 15108 24744
rect 14476 24704 15108 24732
rect 15102 24692 15108 24704
rect 15160 24732 15166 24744
rect 15580 24741 15608 24772
rect 15749 24769 15761 24772
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24800 18567 24803
rect 18598 24800 18604 24812
rect 18555 24772 18604 24800
rect 18555 24769 18567 24772
rect 18509 24763 18567 24769
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 18782 24760 18788 24812
rect 18840 24760 18846 24812
rect 18966 24809 18972 24812
rect 18943 24803 18972 24809
rect 18943 24769 18955 24803
rect 18943 24763 18972 24769
rect 18966 24760 18972 24763
rect 19024 24760 19030 24812
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19352 24800 19380 24840
rect 19291 24772 19380 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 15289 24735 15347 24741
rect 15289 24732 15301 24735
rect 15160 24704 15301 24732
rect 15160 24692 15166 24704
rect 15289 24701 15301 24704
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 15565 24735 15623 24741
rect 15565 24701 15577 24735
rect 15611 24701 15623 24735
rect 15565 24695 15623 24701
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 19076 24732 19104 24760
rect 18463 24704 19104 24732
rect 19168 24732 19196 24763
rect 19426 24760 19432 24812
rect 19484 24760 19490 24812
rect 19536 24800 19564 24840
rect 19610 24828 19616 24880
rect 19668 24868 19674 24880
rect 19886 24868 19892 24880
rect 19668 24840 19892 24868
rect 19668 24828 19674 24840
rect 19886 24828 19892 24840
rect 19944 24868 19950 24880
rect 20165 24871 20223 24877
rect 20165 24868 20177 24871
rect 19944 24840 20177 24868
rect 19944 24828 19950 24840
rect 20165 24837 20177 24840
rect 20211 24837 20223 24871
rect 21266 24868 21272 24880
rect 20165 24831 20223 24837
rect 20364 24840 21272 24868
rect 19536 24772 19932 24800
rect 19168 24704 19564 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 7193 24667 7251 24673
rect 7193 24664 7205 24667
rect 4939 24636 7205 24664
rect 4939 24633 4951 24636
rect 4893 24627 4951 24633
rect 7193 24633 7205 24636
rect 7239 24633 7251 24667
rect 8128 24664 8156 24692
rect 7193 24627 7251 24633
rect 7668 24636 8156 24664
rect 5169 24599 5227 24605
rect 5169 24596 5181 24599
rect 4632 24568 5181 24596
rect 5169 24565 5181 24568
rect 5215 24565 5227 24599
rect 5169 24559 5227 24565
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 6917 24599 6975 24605
rect 6917 24596 6929 24599
rect 6788 24568 6929 24596
rect 6788 24556 6794 24568
rect 6917 24565 6929 24568
rect 6963 24565 6975 24599
rect 6917 24559 6975 24565
rect 7098 24556 7104 24608
rect 7156 24596 7162 24608
rect 7668 24605 7696 24636
rect 12250 24624 12256 24676
rect 12308 24664 12314 24676
rect 13170 24664 13176 24676
rect 12308 24636 13176 24664
rect 12308 24624 12314 24636
rect 13170 24624 13176 24636
rect 13228 24664 13234 24676
rect 13541 24667 13599 24673
rect 13541 24664 13553 24667
rect 13228 24636 13553 24664
rect 13228 24624 13234 24636
rect 13541 24633 13553 24636
rect 13587 24633 13599 24667
rect 13541 24627 13599 24633
rect 18325 24667 18383 24673
rect 18325 24633 18337 24667
rect 18371 24633 18383 24667
rect 18325 24627 18383 24633
rect 18693 24667 18751 24673
rect 18693 24633 18705 24667
rect 18739 24664 18751 24667
rect 19334 24664 19340 24676
rect 18739 24636 19340 24664
rect 18739 24633 18751 24636
rect 18693 24627 18751 24633
rect 7653 24599 7711 24605
rect 7653 24596 7665 24599
rect 7156 24568 7665 24596
rect 7156 24556 7162 24568
rect 7653 24565 7665 24568
rect 7699 24565 7711 24599
rect 7653 24559 7711 24565
rect 7742 24556 7748 24608
rect 7800 24556 7806 24608
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 12529 24599 12587 24605
rect 12529 24596 12541 24599
rect 12492 24568 12541 24596
rect 12492 24556 12498 24568
rect 12529 24565 12541 24568
rect 12575 24565 12587 24599
rect 12529 24559 12587 24565
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13725 24599 13783 24605
rect 13725 24596 13737 24599
rect 13136 24568 13737 24596
rect 13136 24556 13142 24568
rect 13725 24565 13737 24568
rect 13771 24596 13783 24599
rect 13906 24596 13912 24608
rect 13771 24568 13912 24596
rect 13771 24565 13783 24568
rect 13725 24559 13783 24565
rect 13906 24556 13912 24568
rect 13964 24556 13970 24608
rect 18340 24596 18368 24627
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 19536 24673 19564 24704
rect 19794 24692 19800 24744
rect 19852 24692 19858 24744
rect 19904 24732 19932 24772
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 20364 24809 20392 24840
rect 21266 24828 21272 24840
rect 21324 24828 21330 24880
rect 22554 24828 22560 24880
rect 22612 24828 22618 24880
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 20128 24772 20361 24800
rect 20128 24760 20134 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20533 24735 20591 24741
rect 20533 24732 20545 24735
rect 19904 24704 20545 24732
rect 20533 24701 20545 24704
rect 20579 24701 20591 24735
rect 20533 24695 20591 24701
rect 21634 24692 21640 24744
rect 21692 24732 21698 24744
rect 21821 24735 21879 24741
rect 21821 24732 21833 24735
rect 21692 24704 21833 24732
rect 21692 24692 21698 24704
rect 21821 24701 21833 24704
rect 21867 24701 21879 24735
rect 21821 24695 21879 24701
rect 22186 24692 22192 24744
rect 22244 24692 22250 24744
rect 19521 24667 19579 24673
rect 19521 24633 19533 24667
rect 19567 24633 19579 24667
rect 19521 24627 19579 24633
rect 18506 24596 18512 24608
rect 18340 24568 18512 24596
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19705 24599 19763 24605
rect 19705 24596 19717 24599
rect 19208 24568 19717 24596
rect 19208 24556 19214 24568
rect 19705 24565 19717 24568
rect 19751 24565 19763 24599
rect 19705 24559 19763 24565
rect 23290 24556 23296 24608
rect 23348 24596 23354 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 23348 24568 23581 24596
rect 23348 24556 23354 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 1104 24506 26864 24528
rect 1104 24454 4169 24506
rect 4221 24454 4233 24506
rect 4285 24454 4297 24506
rect 4349 24454 4361 24506
rect 4413 24454 4425 24506
rect 4477 24454 10608 24506
rect 10660 24454 10672 24506
rect 10724 24454 10736 24506
rect 10788 24454 10800 24506
rect 10852 24454 10864 24506
rect 10916 24454 17047 24506
rect 17099 24454 17111 24506
rect 17163 24454 17175 24506
rect 17227 24454 17239 24506
rect 17291 24454 17303 24506
rect 17355 24454 23486 24506
rect 23538 24454 23550 24506
rect 23602 24454 23614 24506
rect 23666 24454 23678 24506
rect 23730 24454 23742 24506
rect 23794 24454 26864 24506
rect 1104 24432 26864 24454
rect 3142 24352 3148 24404
rect 3200 24392 3206 24404
rect 3421 24395 3479 24401
rect 3421 24392 3433 24395
rect 3200 24364 3433 24392
rect 3200 24352 3206 24364
rect 3421 24361 3433 24364
rect 3467 24361 3479 24395
rect 3421 24355 3479 24361
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 4525 24395 4583 24401
rect 4525 24392 4537 24395
rect 3936 24364 4537 24392
rect 3936 24352 3942 24364
rect 4525 24361 4537 24364
rect 4571 24361 4583 24395
rect 4525 24355 4583 24361
rect 4709 24395 4767 24401
rect 4709 24361 4721 24395
rect 4755 24392 4767 24395
rect 4798 24392 4804 24404
rect 4755 24364 4804 24392
rect 4755 24361 4767 24364
rect 4709 24355 4767 24361
rect 4062 24284 4068 24336
rect 4120 24284 4126 24336
rect 1394 24216 1400 24268
rect 1452 24216 1458 24268
rect 1765 24259 1823 24265
rect 1765 24225 1777 24259
rect 1811 24256 1823 24259
rect 3694 24256 3700 24268
rect 1811 24228 3700 24256
rect 1811 24225 1823 24228
rect 1765 24219 1823 24225
rect 3694 24216 3700 24228
rect 3752 24216 3758 24268
rect 4522 24256 4528 24268
rect 4264 24228 4528 24256
rect 4264 24200 4292 24228
rect 4522 24216 4528 24228
rect 4580 24256 4586 24268
rect 4724 24256 4752 24355
rect 4798 24352 4804 24364
rect 4856 24392 4862 24404
rect 5534 24392 5540 24404
rect 4856 24364 5540 24392
rect 4856 24352 4862 24364
rect 5534 24352 5540 24364
rect 5592 24352 5598 24404
rect 6273 24395 6331 24401
rect 6273 24361 6285 24395
rect 6319 24392 6331 24395
rect 6546 24392 6552 24404
rect 6319 24364 6552 24392
rect 6319 24361 6331 24364
rect 6273 24355 6331 24361
rect 6546 24352 6552 24364
rect 6604 24352 6610 24404
rect 7006 24401 7012 24404
rect 6963 24395 7012 24401
rect 6963 24361 6975 24395
rect 7009 24361 7012 24395
rect 6963 24355 7012 24361
rect 7006 24352 7012 24355
rect 7064 24352 7070 24404
rect 7101 24395 7159 24401
rect 7101 24361 7113 24395
rect 7147 24392 7159 24395
rect 7650 24392 7656 24404
rect 7147 24364 7656 24392
rect 7147 24361 7159 24364
rect 7101 24355 7159 24361
rect 7650 24352 7656 24364
rect 7708 24352 7714 24404
rect 12894 24352 12900 24404
rect 12952 24392 12958 24404
rect 13173 24395 13231 24401
rect 13173 24392 13185 24395
rect 12952 24364 13185 24392
rect 12952 24352 12958 24364
rect 13173 24361 13185 24364
rect 13219 24361 13231 24395
rect 13173 24355 13231 24361
rect 13262 24352 13268 24404
rect 13320 24392 13326 24404
rect 13357 24395 13415 24401
rect 13357 24392 13369 24395
rect 13320 24364 13369 24392
rect 13320 24352 13326 24364
rect 13357 24361 13369 24364
rect 13403 24392 13415 24395
rect 15930 24392 15936 24404
rect 13403 24364 15936 24392
rect 13403 24361 13415 24364
rect 13357 24355 13415 24361
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 18966 24352 18972 24404
rect 19024 24392 19030 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 19024 24364 19257 24392
rect 19024 24352 19030 24364
rect 19245 24361 19257 24364
rect 19291 24392 19303 24395
rect 19426 24392 19432 24404
rect 19291 24364 19432 24392
rect 19291 24361 19303 24364
rect 19245 24355 19303 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 22281 24395 22339 24401
rect 22281 24361 22293 24395
rect 22327 24392 22339 24395
rect 22554 24392 22560 24404
rect 22327 24364 22560 24392
rect 22327 24361 22339 24364
rect 22281 24355 22339 24361
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 6178 24284 6184 24336
rect 6236 24324 6242 24336
rect 7193 24327 7251 24333
rect 7193 24324 7205 24327
rect 6236 24296 7205 24324
rect 6236 24284 6242 24296
rect 7193 24293 7205 24296
rect 7239 24293 7251 24327
rect 7193 24287 7251 24293
rect 10321 24327 10379 24333
rect 10321 24293 10333 24327
rect 10367 24324 10379 24327
rect 11054 24324 11060 24336
rect 10367 24296 11060 24324
rect 10367 24293 10379 24296
rect 10321 24287 10379 24293
rect 11054 24284 11060 24296
rect 11112 24284 11118 24336
rect 18598 24284 18604 24336
rect 18656 24324 18662 24336
rect 19334 24324 19340 24336
rect 18656 24296 19340 24324
rect 18656 24284 18662 24296
rect 19334 24284 19340 24296
rect 19392 24324 19398 24336
rect 19521 24327 19579 24333
rect 19521 24324 19533 24327
rect 19392 24296 19533 24324
rect 19392 24284 19398 24296
rect 19521 24293 19533 24296
rect 19567 24324 19579 24327
rect 20070 24324 20076 24336
rect 19567 24296 20076 24324
rect 19567 24293 19579 24296
rect 19521 24287 19579 24293
rect 20070 24284 20076 24296
rect 20128 24284 20134 24336
rect 21545 24327 21603 24333
rect 21545 24293 21557 24327
rect 21591 24324 21603 24327
rect 22186 24324 22192 24336
rect 21591 24296 22192 24324
rect 21591 24293 21603 24296
rect 21545 24287 21603 24293
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 7742 24256 7748 24268
rect 4580 24228 4752 24256
rect 6748 24228 7748 24256
rect 4580 24216 4586 24228
rect 2866 24148 2872 24200
rect 2924 24188 2930 24200
rect 3513 24191 3571 24197
rect 3513 24188 3525 24191
rect 2924 24160 3525 24188
rect 2924 24148 2930 24160
rect 3513 24157 3525 24160
rect 3559 24157 3571 24191
rect 3513 24151 3571 24157
rect 3602 24148 3608 24200
rect 3660 24188 3666 24200
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 3660 24160 3985 24188
rect 3660 24148 3666 24160
rect 3973 24157 3985 24160
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4246 24148 4252 24200
rect 4304 24148 4310 24200
rect 4663 24157 4721 24163
rect 2780 24132 2832 24138
rect 4663 24132 4675 24157
rect 3237 24123 3295 24129
rect 3237 24089 3249 24123
rect 3283 24089 3295 24123
rect 3237 24083 3295 24089
rect 2780 24074 2832 24080
rect 3252 24052 3280 24083
rect 4614 24080 4620 24132
rect 4672 24123 4675 24132
rect 4709 24154 4721 24157
rect 4709 24123 4736 24154
rect 4798 24148 4804 24200
rect 4856 24188 4862 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4856 24160 4997 24188
rect 4856 24148 4862 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 5442 24148 5448 24200
rect 5500 24188 5506 24200
rect 6748 24197 6776 24228
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 18506 24216 18512 24268
rect 18564 24256 18570 24268
rect 19613 24259 19671 24265
rect 19613 24256 19625 24259
rect 18564 24228 19625 24256
rect 18564 24216 18570 24228
rect 19613 24225 19625 24228
rect 19659 24225 19671 24259
rect 20438 24256 20444 24268
rect 19613 24219 19671 24225
rect 20088 24228 20444 24256
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 5500 24160 6469 24188
rect 5500 24148 5506 24160
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 6457 24151 6515 24157
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 6825 24191 6883 24197
rect 6825 24157 6837 24191
rect 6871 24188 6883 24191
rect 7098 24188 7104 24200
rect 6871 24160 7104 24188
rect 6871 24157 6883 24160
rect 6825 24151 6883 24157
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24188 7343 24191
rect 7374 24188 7380 24200
rect 7331 24160 7380 24188
rect 7331 24157 7343 24160
rect 7285 24151 7343 24157
rect 7374 24148 7380 24160
rect 7432 24188 7438 24200
rect 8202 24188 8208 24200
rect 7432 24160 8208 24188
rect 7432 24148 7438 24160
rect 8202 24148 8208 24160
rect 8260 24148 8266 24200
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24188 13691 24191
rect 13722 24188 13728 24200
rect 13679 24160 13728 24188
rect 13679 24157 13691 24160
rect 13633 24151 13691 24157
rect 4672 24092 4736 24123
rect 4893 24123 4951 24129
rect 4672 24080 4678 24092
rect 4893 24089 4905 24123
rect 4939 24120 4951 24123
rect 5077 24123 5135 24129
rect 5077 24120 5089 24123
rect 4939 24092 5089 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 5077 24089 5089 24092
rect 5123 24120 5135 24123
rect 10060 24120 10088 24151
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 20088 24197 20116 24228
rect 20438 24216 20444 24228
rect 20496 24256 20502 24268
rect 23290 24256 23296 24268
rect 20496 24228 23296 24256
rect 20496 24216 20502 24228
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19208 24160 19441 24188
rect 19208 24148 19214 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 19981 24191 20039 24197
rect 19981 24188 19993 24191
rect 19751 24160 19993 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 19981 24157 19993 24160
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 5123 24092 10088 24120
rect 10321 24123 10379 24129
rect 5123 24089 5135 24092
rect 5077 24083 5135 24089
rect 10321 24089 10333 24123
rect 10367 24120 10379 24123
rect 10686 24120 10692 24132
rect 10367 24092 10692 24120
rect 10367 24089 10379 24092
rect 10321 24083 10379 24089
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 12986 24080 12992 24132
rect 13044 24080 13050 24132
rect 13170 24080 13176 24132
rect 13228 24129 13234 24132
rect 13228 24123 13247 24129
rect 13235 24089 13247 24123
rect 13228 24083 13247 24089
rect 13228 24080 13234 24083
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 20088 24120 20116 24151
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21324 24160 21373 24188
rect 21324 24148 21330 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24157 21603 24191
rect 21545 24151 21603 24157
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22646 24188 22652 24200
rect 22235 24160 22652 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 19300 24092 20116 24120
rect 19300 24080 19306 24092
rect 20622 24080 20628 24132
rect 20680 24120 20686 24132
rect 21560 24120 21588 24151
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 20680 24092 21588 24120
rect 20680 24080 20686 24092
rect 4246 24052 4252 24064
rect 3252 24024 4252 24052
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 4433 24055 4491 24061
rect 4433 24021 4445 24055
rect 4479 24052 4491 24055
rect 5626 24052 5632 24064
rect 4479 24024 5632 24052
rect 4479 24021 4491 24024
rect 4433 24015 4491 24021
rect 5626 24012 5632 24024
rect 5684 24012 5690 24064
rect 6641 24055 6699 24061
rect 6641 24021 6653 24055
rect 6687 24052 6699 24055
rect 6822 24052 6828 24064
rect 6687 24024 6828 24052
rect 6687 24021 6699 24024
rect 6641 24015 6699 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 10137 24055 10195 24061
rect 10137 24052 10149 24055
rect 10008 24024 10149 24052
rect 10008 24012 10014 24024
rect 10137 24021 10149 24024
rect 10183 24021 10195 24055
rect 10137 24015 10195 24021
rect 13538 24012 13544 24064
rect 13596 24012 13602 24064
rect 21910 24012 21916 24064
rect 21968 24052 21974 24064
rect 22649 24055 22707 24061
rect 22649 24052 22661 24055
rect 21968 24024 22661 24052
rect 21968 24012 21974 24024
rect 22649 24021 22661 24024
rect 22695 24021 22707 24055
rect 22649 24015 22707 24021
rect 1104 23962 26864 23984
rect 1104 23910 4829 23962
rect 4881 23910 4893 23962
rect 4945 23910 4957 23962
rect 5009 23910 5021 23962
rect 5073 23910 5085 23962
rect 5137 23910 11268 23962
rect 11320 23910 11332 23962
rect 11384 23910 11396 23962
rect 11448 23910 11460 23962
rect 11512 23910 11524 23962
rect 11576 23910 17707 23962
rect 17759 23910 17771 23962
rect 17823 23910 17835 23962
rect 17887 23910 17899 23962
rect 17951 23910 17963 23962
rect 18015 23910 24146 23962
rect 24198 23910 24210 23962
rect 24262 23910 24274 23962
rect 24326 23910 24338 23962
rect 24390 23910 24402 23962
rect 24454 23910 26864 23962
rect 1104 23888 26864 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 1627 23820 2268 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 2240 23789 2268 23820
rect 2774 23808 2780 23860
rect 2832 23808 2838 23860
rect 3970 23808 3976 23860
rect 4028 23848 4034 23860
rect 4157 23851 4215 23857
rect 4157 23848 4169 23851
rect 4028 23820 4169 23848
rect 4028 23808 4034 23820
rect 4157 23817 4169 23820
rect 4203 23817 4215 23851
rect 4157 23811 4215 23817
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 8202 23857 8208 23860
rect 8159 23851 8208 23857
rect 5592 23820 7880 23848
rect 5592 23808 5598 23820
rect 2225 23783 2283 23789
rect 2225 23749 2237 23783
rect 2271 23749 2283 23783
rect 4246 23780 4252 23792
rect 2225 23743 2283 23749
rect 3896 23752 4252 23780
rect 934 23672 940 23724
rect 992 23712 998 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 992 23684 1409 23712
rect 992 23672 998 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 2866 23672 2872 23724
rect 2924 23672 2930 23724
rect 3896 23721 3924 23752
rect 4246 23740 4252 23752
rect 4304 23740 4310 23792
rect 7098 23740 7104 23792
rect 7156 23740 7162 23792
rect 7852 23780 7880 23820
rect 8159 23817 8171 23851
rect 8205 23817 8208 23851
rect 8159 23811 8208 23817
rect 8202 23808 8208 23811
rect 8260 23808 8266 23860
rect 10226 23848 10232 23860
rect 9416 23820 10232 23848
rect 9306 23780 9312 23792
rect 7852 23752 9312 23780
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23681 3939 23715
rect 3881 23675 3939 23681
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23712 4031 23715
rect 4614 23712 4620 23724
rect 4019 23684 4620 23712
rect 4019 23681 4031 23684
rect 3973 23675 4031 23681
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6365 23715 6423 23721
rect 6365 23712 6377 23715
rect 6328 23684 6377 23712
rect 6328 23672 6334 23684
rect 6365 23681 6377 23684
rect 6411 23712 6423 23715
rect 6638 23712 6644 23724
rect 6411 23684 6644 23712
rect 6411 23681 6423 23684
rect 6365 23675 6423 23681
rect 6638 23672 6644 23684
rect 6696 23672 6702 23724
rect 6730 23672 6736 23724
rect 6788 23672 6794 23724
rect 9214 23672 9220 23724
rect 9272 23672 9278 23724
rect 9416 23721 9444 23820
rect 10226 23808 10232 23820
rect 10284 23808 10290 23860
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 13541 23851 13599 23857
rect 10560 23820 12434 23848
rect 10560 23808 10566 23820
rect 12406 23780 12434 23820
rect 13541 23817 13553 23851
rect 13587 23848 13599 23851
rect 13814 23848 13820 23860
rect 13587 23820 13820 23848
rect 13587 23817 13599 23820
rect 13541 23811 13599 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 19794 23808 19800 23860
rect 19852 23808 19858 23860
rect 21376 23820 22094 23848
rect 13078 23780 13084 23792
rect 12406 23752 13084 23780
rect 13078 23740 13084 23752
rect 13136 23740 13142 23792
rect 14645 23783 14703 23789
rect 14645 23780 14657 23783
rect 13924 23752 14657 23780
rect 10318 23721 10324 23724
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23681 9459 23715
rect 9401 23675 9459 23681
rect 10296 23715 10324 23721
rect 10296 23681 10308 23715
rect 10296 23675 10324 23681
rect 10318 23672 10324 23675
rect 10376 23672 10382 23724
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23681 10471 23715
rect 10413 23675 10471 23681
rect 11333 23715 11391 23721
rect 11333 23681 11345 23715
rect 11379 23712 11391 23715
rect 11698 23712 11704 23724
rect 11379 23684 11704 23712
rect 11379 23681 11391 23684
rect 11333 23675 11391 23681
rect 4154 23604 4160 23656
rect 4212 23604 4218 23656
rect 4706 23604 4712 23656
rect 4764 23644 4770 23656
rect 9766 23644 9772 23656
rect 4764 23616 9772 23644
rect 4764 23604 4770 23616
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 9950 23604 9956 23656
rect 10008 23644 10014 23656
rect 10137 23647 10195 23653
rect 10137 23644 10149 23647
rect 10008 23616 10149 23644
rect 10008 23604 10014 23616
rect 10137 23613 10149 23616
rect 10183 23613 10195 23647
rect 10428 23644 10456 23675
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 12676 23684 13461 23712
rect 12676 23672 12682 23684
rect 13449 23681 13461 23684
rect 13495 23712 13507 23715
rect 13538 23712 13544 23724
rect 13495 23684 13544 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13814 23712 13820 23724
rect 13679 23684 13820 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 13814 23672 13820 23684
rect 13872 23672 13878 23724
rect 13924 23721 13952 23752
rect 14645 23749 14657 23752
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 18230 23740 18236 23792
rect 18288 23780 18294 23792
rect 19150 23780 19156 23792
rect 18288 23752 19156 23780
rect 18288 23740 18294 23752
rect 19150 23740 19156 23752
rect 19208 23780 19214 23792
rect 19245 23783 19303 23789
rect 19245 23780 19257 23783
rect 19208 23752 19257 23780
rect 19208 23740 19214 23752
rect 19245 23749 19257 23752
rect 19291 23749 19303 23783
rect 19245 23743 19303 23749
rect 19475 23749 19533 23755
rect 19475 23746 19487 23749
rect 13909 23715 13967 23721
rect 13909 23681 13921 23715
rect 13955 23681 13967 23715
rect 13909 23675 13967 23681
rect 14369 23715 14427 23721
rect 14369 23681 14381 23715
rect 14415 23712 14427 23715
rect 14826 23712 14832 23724
rect 14415 23684 14832 23712
rect 14415 23681 14427 23684
rect 14369 23675 14427 23681
rect 14826 23672 14832 23684
rect 14884 23712 14890 23724
rect 16393 23715 16451 23721
rect 16393 23712 16405 23715
rect 14884 23684 16405 23712
rect 14884 23672 14890 23684
rect 16393 23681 16405 23684
rect 16439 23681 16451 23715
rect 19334 23712 19340 23724
rect 16393 23675 16451 23681
rect 19260 23684 19340 23712
rect 10594 23644 10600 23656
rect 10428 23616 10600 23644
rect 10137 23607 10195 23613
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 11149 23647 11207 23653
rect 11149 23613 11161 23647
rect 11195 23613 11207 23647
rect 11149 23607 11207 23613
rect 4172 23576 4200 23604
rect 5258 23576 5264 23588
rect 4172 23548 5264 23576
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 9401 23579 9459 23585
rect 9401 23545 9413 23579
rect 9447 23576 9459 23579
rect 9447 23548 9812 23576
rect 9447 23545 9459 23548
rect 9401 23539 9459 23545
rect 2501 23511 2559 23517
rect 2501 23477 2513 23511
rect 2547 23508 2559 23511
rect 2774 23508 2780 23520
rect 2547 23480 2780 23508
rect 2547 23477 2559 23480
rect 2501 23471 2559 23477
rect 2774 23468 2780 23480
rect 2832 23468 2838 23520
rect 9493 23511 9551 23517
rect 9493 23477 9505 23511
rect 9539 23508 9551 23511
rect 9674 23508 9680 23520
rect 9539 23480 9680 23508
rect 9539 23477 9551 23480
rect 9493 23471 9551 23477
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 9784 23508 9812 23548
rect 10686 23536 10692 23588
rect 10744 23576 10750 23588
rect 11164 23576 11192 23607
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 10744 23548 11100 23576
rect 11164 23548 18920 23576
rect 10744 23536 10750 23548
rect 10962 23508 10968 23520
rect 9784 23480 10968 23508
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 11072 23508 11100 23548
rect 12066 23508 12072 23520
rect 11072 23480 12072 23508
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 13814 23468 13820 23520
rect 13872 23468 13878 23520
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 14461 23511 14519 23517
rect 14461 23508 14473 23511
rect 14424 23480 14473 23508
rect 14424 23468 14430 23480
rect 14461 23477 14473 23480
rect 14507 23477 14519 23511
rect 14461 23471 14519 23477
rect 16298 23468 16304 23520
rect 16356 23468 16362 23520
rect 18892 23508 18920 23548
rect 19260 23508 19288 23684
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 19465 23715 19487 23746
rect 19521 23715 19533 23749
rect 19465 23712 19533 23715
rect 19705 23715 19763 23721
rect 19705 23712 19717 23715
rect 19465 23684 19717 23712
rect 19705 23681 19717 23684
rect 19751 23712 19763 23715
rect 19886 23712 19892 23724
rect 19751 23684 19892 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 20898 23672 20904 23724
rect 20956 23712 20962 23724
rect 21376 23721 21404 23820
rect 21637 23783 21695 23789
rect 21637 23749 21649 23783
rect 21683 23780 21695 23783
rect 21910 23780 21916 23792
rect 21683 23752 21916 23780
rect 21683 23749 21695 23752
rect 21637 23743 21695 23749
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22066 23780 22094 23820
rect 22186 23808 22192 23860
rect 22244 23848 22250 23860
rect 22465 23851 22523 23857
rect 22465 23848 22477 23851
rect 22244 23820 22477 23848
rect 22244 23808 22250 23820
rect 22465 23817 22477 23820
rect 22511 23817 22523 23851
rect 22465 23811 22523 23817
rect 22066 23752 22600 23780
rect 21361 23715 21419 23721
rect 21361 23712 21373 23715
rect 20956 23684 21373 23712
rect 20956 23672 20962 23684
rect 21361 23681 21373 23684
rect 21407 23681 21419 23715
rect 21361 23675 21419 23681
rect 21450 23672 21456 23724
rect 21508 23672 21514 23724
rect 21542 23672 21548 23724
rect 21600 23712 21606 23724
rect 22572 23721 22600 23752
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21600 23684 21833 23712
rect 21600 23672 21606 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 20622 23644 20628 23656
rect 19628 23616 20628 23644
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 19628 23585 19656 23616
rect 20622 23604 20628 23616
rect 20680 23644 20686 23656
rect 22020 23644 22048 23675
rect 20680 23616 22048 23644
rect 20680 23604 20686 23616
rect 19613 23579 19671 23585
rect 19613 23576 19625 23579
rect 19392 23548 19625 23576
rect 19392 23536 19398 23548
rect 19613 23545 19625 23548
rect 19659 23545 19671 23579
rect 19613 23539 19671 23545
rect 21637 23579 21695 23585
rect 21637 23545 21649 23579
rect 21683 23576 21695 23579
rect 22296 23576 22324 23675
rect 22646 23672 22652 23724
rect 22704 23672 22710 23724
rect 21683 23548 22324 23576
rect 21683 23545 21695 23548
rect 21637 23539 21695 23545
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 18892 23480 19441 23508
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 19429 23471 19487 23477
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22189 23511 22247 23517
rect 22189 23508 22201 23511
rect 22152 23480 22201 23508
rect 22152 23468 22158 23480
rect 22189 23477 22201 23480
rect 22235 23477 22247 23511
rect 22189 23471 22247 23477
rect 22278 23468 22284 23520
rect 22336 23468 22342 23520
rect 22646 23468 22652 23520
rect 22704 23508 22710 23520
rect 22741 23511 22799 23517
rect 22741 23508 22753 23511
rect 22704 23480 22753 23508
rect 22704 23468 22710 23480
rect 22741 23477 22753 23480
rect 22787 23477 22799 23511
rect 22741 23471 22799 23477
rect 1104 23418 26864 23440
rect 1104 23366 4169 23418
rect 4221 23366 4233 23418
rect 4285 23366 4297 23418
rect 4349 23366 4361 23418
rect 4413 23366 4425 23418
rect 4477 23366 10608 23418
rect 10660 23366 10672 23418
rect 10724 23366 10736 23418
rect 10788 23366 10800 23418
rect 10852 23366 10864 23418
rect 10916 23366 17047 23418
rect 17099 23366 17111 23418
rect 17163 23366 17175 23418
rect 17227 23366 17239 23418
rect 17291 23366 17303 23418
rect 17355 23366 23486 23418
rect 23538 23366 23550 23418
rect 23602 23366 23614 23418
rect 23666 23366 23678 23418
rect 23730 23366 23742 23418
rect 23794 23366 26864 23418
rect 1104 23344 26864 23366
rect 7098 23264 7104 23316
rect 7156 23264 7162 23316
rect 8573 23307 8631 23313
rect 8573 23273 8585 23307
rect 8619 23304 8631 23307
rect 9122 23304 9128 23316
rect 8619 23276 9128 23304
rect 8619 23273 8631 23276
rect 8573 23267 8631 23273
rect 9122 23264 9128 23276
rect 9180 23264 9186 23316
rect 9398 23264 9404 23316
rect 9456 23304 9462 23316
rect 9456 23276 10180 23304
rect 9456 23264 9462 23276
rect 8110 23196 8116 23248
rect 8168 23236 8174 23248
rect 8938 23236 8944 23248
rect 8168 23208 8944 23236
rect 8168 23196 8174 23208
rect 8938 23196 8944 23208
rect 8996 23196 9002 23248
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 3053 23171 3111 23177
rect 3053 23168 3065 23171
rect 2924 23140 3065 23168
rect 2924 23128 2930 23140
rect 3053 23137 3065 23140
rect 3099 23168 3111 23171
rect 3099 23140 6408 23168
rect 3099 23137 3111 23140
rect 3053 23131 3111 23137
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 3234 23100 3240 23112
rect 2832 23072 3240 23100
rect 2832 23060 2838 23072
rect 3234 23060 3240 23072
rect 3292 23100 3298 23112
rect 6178 23100 6184 23112
rect 3292 23072 6184 23100
rect 3292 23060 3298 23072
rect 6178 23060 6184 23072
rect 6236 23100 6242 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 6236 23072 6285 23100
rect 6236 23060 6242 23072
rect 6273 23069 6285 23072
rect 6319 23069 6331 23103
rect 6380 23100 6408 23140
rect 6730 23128 6736 23180
rect 6788 23168 6794 23180
rect 9030 23168 9036 23180
rect 6788 23140 9036 23168
rect 6788 23128 6794 23140
rect 9030 23128 9036 23140
rect 9088 23128 9094 23180
rect 9582 23128 9588 23180
rect 9640 23128 9646 23180
rect 9858 23128 9864 23180
rect 9916 23128 9922 23180
rect 10152 23177 10180 23276
rect 10502 23264 10508 23316
rect 10560 23304 10566 23316
rect 11701 23307 11759 23313
rect 10560 23276 10824 23304
rect 10560 23264 10566 23276
rect 10137 23171 10195 23177
rect 10137 23137 10149 23171
rect 10183 23168 10195 23171
rect 10183 23140 10456 23168
rect 10183 23137 10195 23140
rect 10137 23131 10195 23137
rect 7009 23103 7067 23109
rect 7009 23100 7021 23103
rect 6380 23072 7021 23100
rect 6273 23063 6331 23069
rect 7009 23069 7021 23072
rect 7055 23100 7067 23103
rect 7098 23100 7104 23112
rect 7055 23072 7104 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23100 8263 23103
rect 8386 23100 8392 23112
rect 8251 23072 8392 23100
rect 8251 23069 8263 23072
rect 8205 23063 8263 23069
rect 8386 23060 8392 23072
rect 8444 23060 8450 23112
rect 9766 23109 9772 23112
rect 9744 23103 9772 23109
rect 9744 23069 9756 23103
rect 9744 23063 9772 23069
rect 9766 23060 9772 23063
rect 9824 23060 9830 23112
rect 10428 23100 10456 23140
rect 10502 23128 10508 23180
rect 10560 23168 10566 23180
rect 10796 23177 10824 23276
rect 11701 23273 11713 23307
rect 11747 23304 11759 23307
rect 12434 23304 12440 23316
rect 11747 23276 12440 23304
rect 11747 23273 11759 23276
rect 11701 23267 11759 23273
rect 12434 23264 12440 23276
rect 12492 23264 12498 23316
rect 12802 23264 12808 23316
rect 12860 23304 12866 23316
rect 12897 23307 12955 23313
rect 12897 23304 12909 23307
rect 12860 23276 12909 23304
rect 12860 23264 12866 23276
rect 12897 23273 12909 23276
rect 12943 23273 12955 23307
rect 12897 23267 12955 23273
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 15654 23304 15660 23316
rect 15519 23276 15660 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23304 18475 23307
rect 19702 23304 19708 23316
rect 18463 23276 19708 23304
rect 18463 23273 18475 23276
rect 18417 23267 18475 23273
rect 19702 23264 19708 23276
rect 19760 23264 19766 23316
rect 19886 23264 19892 23316
rect 19944 23264 19950 23316
rect 20070 23264 20076 23316
rect 20128 23264 20134 23316
rect 20898 23264 20904 23316
rect 20956 23264 20962 23316
rect 22094 23304 22100 23316
rect 21284 23276 22100 23304
rect 11790 23196 11796 23248
rect 11848 23236 11854 23248
rect 12345 23239 12403 23245
rect 12345 23236 12357 23239
rect 11848 23208 12357 23236
rect 11848 23196 11854 23208
rect 12345 23205 12357 23208
rect 12391 23205 12403 23239
rect 12345 23199 12403 23205
rect 12986 23196 12992 23248
rect 13044 23236 13050 23248
rect 13357 23239 13415 23245
rect 13357 23236 13369 23239
rect 13044 23208 13369 23236
rect 13044 23196 13050 23208
rect 13357 23205 13369 23208
rect 13403 23205 13415 23239
rect 19334 23236 19340 23248
rect 13357 23199 13415 23205
rect 18892 23208 19340 23236
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 10560 23140 10609 23168
rect 10560 23128 10566 23140
rect 10597 23137 10609 23140
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 10781 23171 10839 23177
rect 10781 23137 10793 23171
rect 10827 23137 10839 23171
rect 10781 23131 10839 23137
rect 11333 23171 11391 23177
rect 11333 23137 11345 23171
rect 11379 23168 11391 23171
rect 12158 23168 12164 23180
rect 11379 23140 12164 23168
rect 11379 23137 11391 23140
rect 11333 23131 11391 23137
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 13265 23171 13323 23177
rect 12360 23140 12756 23168
rect 10686 23100 10692 23112
rect 10428 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 11054 23060 11060 23112
rect 11112 23060 11118 23112
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 11422 23060 11428 23112
rect 11480 23060 11486 23112
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 12360 23109 12388 23140
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 11940 23072 12081 23100
rect 11940 23060 11946 23072
rect 12069 23069 12081 23072
rect 12115 23100 12127 23103
rect 12345 23103 12403 23109
rect 12345 23100 12357 23103
rect 12115 23072 12357 23100
rect 12115 23069 12127 23072
rect 12069 23063 12127 23069
rect 12345 23069 12357 23072
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12728 23100 12756 23140
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 14182 23168 14188 23180
rect 13311 23140 14188 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 16666 23128 16672 23180
rect 16724 23168 16730 23180
rect 17221 23171 17279 23177
rect 17221 23168 17233 23171
rect 16724 23140 17233 23168
rect 16724 23128 16730 23140
rect 17221 23137 17233 23140
rect 17267 23137 17279 23171
rect 17221 23131 17279 23137
rect 13633 23103 13691 23109
rect 12728 23072 13308 23100
rect 5994 22992 6000 23044
rect 6052 22992 6058 23044
rect 8018 22992 8024 23044
rect 8076 23032 8082 23044
rect 8573 23035 8631 23041
rect 8573 23032 8585 23035
rect 8076 23004 8585 23032
rect 8076 22992 8082 23004
rect 8573 23001 8585 23004
rect 8619 23001 8631 23035
rect 8573 22995 8631 23001
rect 10873 23035 10931 23041
rect 10873 23001 10885 23035
rect 10919 23032 10931 23035
rect 11716 23032 11744 23060
rect 13280 23044 13308 23072
rect 13633 23069 13645 23103
rect 13679 23100 13691 23103
rect 13814 23100 13820 23112
rect 13679 23072 13820 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 16850 23060 16856 23112
rect 16908 23060 16914 23112
rect 18322 23060 18328 23112
rect 18380 23060 18386 23112
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 18892 23100 18920 23208
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 19812 23140 21128 23168
rect 18831 23072 18920 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 19058 23060 19064 23112
rect 19116 23060 19122 23112
rect 19242 23060 19248 23112
rect 19300 23060 19306 23112
rect 19518 23060 19524 23112
rect 19576 23060 19582 23112
rect 19702 23109 19708 23112
rect 19659 23103 19708 23109
rect 19659 23069 19671 23103
rect 19705 23069 19708 23103
rect 19659 23063 19708 23069
rect 19702 23060 19708 23063
rect 19760 23060 19766 23112
rect 10919 23004 11744 23032
rect 12529 23035 12587 23041
rect 10919 23001 10931 23004
rect 10873 22995 10931 23001
rect 12529 23001 12541 23035
rect 12575 23032 12587 23035
rect 12575 23004 13032 23032
rect 12575 23001 12587 23004
rect 12529 22995 12587 23001
rect 8757 22967 8815 22973
rect 8757 22933 8769 22967
rect 8803 22964 8815 22967
rect 8846 22964 8852 22976
rect 8803 22936 8852 22964
rect 8803 22933 8815 22936
rect 8757 22927 8815 22933
rect 8846 22924 8852 22936
rect 8904 22924 8910 22976
rect 8941 22967 8999 22973
rect 8941 22933 8953 22967
rect 8987 22964 8999 22967
rect 10226 22964 10232 22976
rect 8987 22936 10232 22964
rect 8987 22933 8999 22936
rect 8941 22927 8999 22933
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 11517 22967 11575 22973
rect 11517 22933 11529 22967
rect 11563 22964 11575 22967
rect 11606 22964 11612 22976
rect 11563 22936 11612 22964
rect 11563 22933 11575 22936
rect 11517 22927 11575 22933
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22964 11759 22967
rect 12066 22964 12072 22976
rect 11747 22936 12072 22964
rect 11747 22933 11759 22936
rect 11701 22927 11759 22933
rect 12066 22924 12072 22936
rect 12124 22964 12130 22976
rect 12544 22964 12572 22995
rect 12124 22936 12572 22964
rect 12124 22924 12130 22936
rect 12710 22924 12716 22976
rect 12768 22924 12774 22976
rect 12894 22924 12900 22976
rect 12952 22924 12958 22976
rect 13004 22964 13032 23004
rect 13262 22992 13268 23044
rect 13320 23032 13326 23044
rect 13357 23035 13415 23041
rect 13357 23032 13369 23035
rect 13320 23004 13369 23032
rect 13320 22992 13326 23004
rect 13357 23001 13369 23004
rect 13403 23001 13415 23035
rect 13357 22995 13415 23001
rect 16298 22992 16304 23044
rect 16356 22992 16362 23044
rect 18601 23035 18659 23041
rect 18601 23001 18613 23035
rect 18647 23032 18659 23035
rect 19429 23035 19487 23041
rect 19429 23032 19441 23035
rect 18647 23004 19441 23032
rect 18647 23001 18659 23004
rect 18601 22995 18659 23001
rect 19429 23001 19441 23004
rect 19475 23001 19487 23035
rect 19536 23032 19564 23060
rect 19812 23032 19840 23140
rect 20438 23060 20444 23112
rect 20496 23100 20502 23112
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20496 23072 21005 23100
rect 20496 23060 20502 23072
rect 20993 23069 21005 23072
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 19536 23004 19840 23032
rect 19429 22995 19487 23001
rect 19886 22992 19892 23044
rect 19944 23032 19950 23044
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 19944 23004 20269 23032
rect 19944 22992 19950 23004
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20530 23032 20536 23044
rect 20588 23041 20594 23044
rect 20588 23035 20609 23041
rect 20257 22995 20315 23001
rect 20456 23004 20536 23032
rect 13446 22964 13452 22976
rect 13004 22936 13452 22964
rect 13446 22924 13452 22936
rect 13504 22964 13510 22976
rect 13541 22967 13599 22973
rect 13541 22964 13553 22967
rect 13504 22936 13553 22964
rect 13504 22924 13510 22936
rect 13541 22933 13553 22936
rect 13587 22933 13599 22967
rect 13541 22927 13599 22933
rect 18969 22967 19027 22973
rect 18969 22933 18981 22967
rect 19015 22964 19027 22967
rect 19610 22964 19616 22976
rect 19015 22936 19616 22964
rect 19015 22933 19027 22936
rect 18969 22927 19027 22933
rect 19610 22924 19616 22936
rect 19668 22924 19674 22976
rect 19794 22924 19800 22976
rect 19852 22924 19858 22976
rect 20057 22967 20115 22973
rect 20057 22933 20069 22967
rect 20103 22964 20115 22967
rect 20456 22964 20484 23004
rect 20530 22992 20536 23004
rect 20597 23001 20609 23035
rect 20588 22995 20609 23001
rect 20588 22992 20594 22995
rect 20714 22992 20720 23044
rect 20772 22992 20778 23044
rect 21100 23032 21128 23140
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23100 21235 23103
rect 21284 23100 21312 23276
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 21913 23171 21971 23177
rect 21913 23137 21925 23171
rect 21959 23168 21971 23171
rect 22278 23168 22284 23180
rect 21959 23140 22284 23168
rect 21959 23137 21971 23140
rect 21913 23131 21971 23137
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 21223 23072 21312 23100
rect 21223 23069 21235 23072
rect 21177 23063 21235 23069
rect 21358 23060 21364 23112
rect 21416 23060 21422 23112
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21266 23032 21272 23044
rect 21100 23004 21272 23032
rect 21266 22992 21272 23004
rect 21324 22992 21330 23044
rect 21376 23004 22232 23032
rect 20103 22936 20484 22964
rect 20103 22933 20115 22936
rect 20057 22927 20115 22933
rect 20806 22924 20812 22976
rect 20864 22964 20870 22976
rect 21376 22964 21404 23004
rect 20864 22936 21404 22964
rect 21545 22967 21603 22973
rect 20864 22924 20870 22936
rect 21545 22933 21557 22967
rect 21591 22964 21603 22967
rect 22094 22964 22100 22976
rect 21591 22936 22100 22964
rect 21591 22933 21603 22936
rect 21545 22927 21603 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22204 22964 22232 23004
rect 22646 22992 22652 23044
rect 22704 22992 22710 23044
rect 23385 22967 23443 22973
rect 23385 22964 23397 22967
rect 22204 22936 23397 22964
rect 23385 22933 23397 22936
rect 23431 22933 23443 22967
rect 23385 22927 23443 22933
rect 1104 22874 26864 22896
rect 1104 22822 4829 22874
rect 4881 22822 4893 22874
rect 4945 22822 4957 22874
rect 5009 22822 5021 22874
rect 5073 22822 5085 22874
rect 5137 22822 11268 22874
rect 11320 22822 11332 22874
rect 11384 22822 11396 22874
rect 11448 22822 11460 22874
rect 11512 22822 11524 22874
rect 11576 22822 17707 22874
rect 17759 22822 17771 22874
rect 17823 22822 17835 22874
rect 17887 22822 17899 22874
rect 17951 22822 17963 22874
rect 18015 22822 24146 22874
rect 24198 22822 24210 22874
rect 24262 22822 24274 22874
rect 24326 22822 24338 22874
rect 24390 22822 24402 22874
rect 24454 22822 26864 22874
rect 1104 22800 26864 22822
rect 6546 22720 6552 22772
rect 6604 22760 6610 22772
rect 9585 22763 9643 22769
rect 6604 22732 9444 22760
rect 6604 22720 6610 22732
rect 8202 22652 8208 22704
rect 8260 22692 8266 22704
rect 8757 22695 8815 22701
rect 8757 22692 8769 22695
rect 8260 22664 8769 22692
rect 8260 22652 8266 22664
rect 8757 22661 8769 22664
rect 8803 22661 8815 22695
rect 8757 22655 8815 22661
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 8846 22584 8852 22636
rect 8904 22624 8910 22636
rect 9416 22633 9444 22732
rect 9585 22729 9597 22763
rect 9631 22760 9643 22763
rect 9631 22732 11008 22760
rect 9631 22729 9643 22732
rect 9585 22723 9643 22729
rect 10980 22692 11008 22732
rect 11514 22720 11520 22772
rect 11572 22760 11578 22772
rect 11882 22760 11888 22772
rect 11572 22732 11888 22760
rect 11572 22720 11578 22732
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 11974 22720 11980 22772
rect 12032 22760 12038 22772
rect 12805 22763 12863 22769
rect 12032 22732 12572 22760
rect 12032 22720 12038 22732
rect 12434 22692 12440 22704
rect 10980 22664 11744 22692
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8904 22596 9137 22624
rect 8904 22584 8910 22596
rect 9125 22593 9137 22596
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9674 22584 9680 22636
rect 9732 22584 9738 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22593 10011 22627
rect 9953 22587 10011 22593
rect 9214 22516 9220 22568
rect 9272 22516 9278 22568
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22556 9367 22559
rect 9490 22556 9496 22568
rect 9355 22528 9496 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 8941 22491 8999 22497
rect 8941 22457 8953 22491
rect 8987 22488 8999 22491
rect 8987 22460 9720 22488
rect 8987 22457 8999 22460
rect 8941 22451 8999 22457
rect 8757 22423 8815 22429
rect 8757 22389 8769 22423
rect 8803 22420 8815 22423
rect 9122 22420 9128 22432
rect 8803 22392 9128 22420
rect 8803 22389 8815 22392
rect 8757 22383 8815 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 9692 22429 9720 22460
rect 9858 22448 9864 22500
rect 9916 22488 9922 22500
rect 9968 22488 9996 22587
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10781 22627 10839 22633
rect 10781 22624 10793 22627
rect 10192 22596 10793 22624
rect 10192 22584 10198 22596
rect 10781 22593 10793 22596
rect 10827 22593 10839 22627
rect 10781 22587 10839 22593
rect 10962 22584 10968 22636
rect 11020 22584 11026 22636
rect 11716 22633 11744 22664
rect 12084 22664 12440 22692
rect 11241 22627 11299 22633
rect 11241 22593 11253 22627
rect 11287 22593 11299 22627
rect 11241 22587 11299 22593
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11054 22516 11060 22568
rect 11112 22516 11118 22568
rect 11256 22556 11284 22587
rect 11790 22584 11796 22636
rect 11848 22584 11854 22636
rect 12084 22633 12112 22664
rect 12434 22652 12440 22664
rect 12492 22652 12498 22704
rect 12544 22692 12572 22732
rect 12805 22729 12817 22763
rect 12851 22760 12863 22763
rect 13446 22760 13452 22772
rect 12851 22732 13452 22760
rect 12851 22729 12863 22732
rect 12805 22723 12863 22729
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 15194 22720 15200 22772
rect 15252 22769 15258 22772
rect 15252 22763 15301 22769
rect 15252 22729 15255 22763
rect 15289 22729 15301 22763
rect 15252 22723 15301 22729
rect 15252 22720 15258 22723
rect 16942 22720 16948 22772
rect 17000 22760 17006 22772
rect 17000 22732 20576 22760
rect 17000 22720 17006 22732
rect 12544 22664 13032 22692
rect 12544 22633 12572 22664
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12529 22627 12587 22633
rect 12391 22596 12480 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12452 22568 12480 22596
rect 12529 22593 12541 22627
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22624 12679 22627
rect 12894 22624 12900 22636
rect 12667 22596 12900 22624
rect 12667 22593 12679 22596
rect 12621 22587 12679 22593
rect 12250 22556 12256 22568
rect 11256 22528 12256 22556
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 12636 22556 12664 22587
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13004 22624 13032 22664
rect 14366 22652 14372 22704
rect 14424 22652 14430 22704
rect 17954 22652 17960 22704
rect 18012 22652 18018 22704
rect 19978 22692 19984 22704
rect 19826 22664 19984 22692
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 20548 22692 20576 22732
rect 21634 22692 21640 22704
rect 20548 22664 21640 22692
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 13004 22596 13093 22624
rect 13081 22593 13093 22596
rect 13127 22593 13139 22627
rect 13081 22587 13139 22593
rect 12492 22528 12664 22556
rect 13096 22556 13124 22587
rect 13354 22584 13360 22636
rect 13412 22624 13418 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 13412 22596 13461 22624
rect 13412 22584 13418 22596
rect 13449 22593 13461 22596
rect 13495 22593 13507 22627
rect 13449 22587 13507 22593
rect 13814 22584 13820 22636
rect 13872 22584 13878 22636
rect 15838 22584 15844 22636
rect 15896 22584 15902 22636
rect 16666 22584 16672 22636
rect 16724 22584 16730 22636
rect 20548 22633 20576 22664
rect 21634 22652 21640 22664
rect 21692 22692 21698 22704
rect 21692 22664 21864 22692
rect 21692 22652 21698 22664
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20622 22584 20628 22636
rect 20680 22584 20686 22636
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 21836 22633 21864 22664
rect 22094 22652 22100 22704
rect 22152 22652 22158 22704
rect 22646 22652 22652 22704
rect 22704 22652 22710 22704
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22624 21143 22627
rect 21821 22627 21879 22633
rect 21131 22596 21680 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 21652 22568 21680 22596
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 14182 22556 14188 22568
rect 13096 22528 14188 22556
rect 12492 22516 12498 22528
rect 14182 22516 14188 22528
rect 14240 22516 14246 22568
rect 16117 22559 16175 22565
rect 16117 22525 16129 22559
rect 16163 22556 16175 22559
rect 16574 22556 16580 22568
rect 16163 22528 16580 22556
rect 16163 22525 16175 22528
rect 16117 22519 16175 22525
rect 16574 22516 16580 22528
rect 16632 22516 16638 22568
rect 16945 22559 17003 22565
rect 16945 22556 16957 22559
rect 16776 22528 16957 22556
rect 9916 22460 9996 22488
rect 10873 22491 10931 22497
rect 9916 22448 9922 22460
rect 10873 22457 10885 22491
rect 10919 22488 10931 22491
rect 12986 22488 12992 22500
rect 10919 22460 12992 22488
rect 10919 22457 10931 22460
rect 10873 22451 10931 22457
rect 12986 22448 12992 22460
rect 13044 22448 13050 22500
rect 16776 22432 16804 22528
rect 16945 22525 16957 22528
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 18693 22559 18751 22565
rect 18693 22556 18705 22559
rect 18656 22528 18705 22556
rect 18656 22516 18662 22528
rect 18693 22525 18705 22528
rect 18739 22525 18751 22559
rect 18693 22519 18751 22525
rect 18782 22516 18788 22568
rect 18840 22556 18846 22568
rect 19702 22556 19708 22568
rect 18840 22528 19708 22556
rect 18840 22516 18846 22528
rect 19702 22516 19708 22528
rect 19760 22516 19766 22568
rect 19794 22516 19800 22568
rect 19852 22556 19858 22568
rect 20257 22559 20315 22565
rect 20257 22556 20269 22559
rect 19852 22528 20269 22556
rect 19852 22516 19858 22528
rect 20257 22525 20269 22528
rect 20303 22525 20315 22559
rect 20257 22519 20315 22525
rect 20993 22559 21051 22565
rect 20993 22525 21005 22559
rect 21039 22525 21051 22559
rect 20993 22519 21051 22525
rect 21453 22559 21511 22565
rect 21453 22525 21465 22559
rect 21499 22556 21511 22559
rect 21542 22556 21548 22568
rect 21499 22528 21548 22556
rect 21499 22525 21511 22528
rect 21453 22519 21511 22525
rect 20530 22448 20536 22500
rect 20588 22488 20594 22500
rect 21008 22488 21036 22519
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 21692 22528 23857 22556
rect 21692 22516 21698 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 20588 22460 21036 22488
rect 20588 22448 20594 22460
rect 9677 22423 9735 22429
rect 9677 22389 9689 22423
rect 9723 22389 9735 22423
rect 9677 22383 9735 22389
rect 10042 22380 10048 22432
rect 10100 22420 10106 22432
rect 10137 22423 10195 22429
rect 10137 22420 10149 22423
rect 10100 22392 10149 22420
rect 10100 22380 10106 22392
rect 10137 22389 10149 22392
rect 10183 22389 10195 22423
rect 10137 22383 10195 22389
rect 10410 22380 10416 22432
rect 10468 22420 10474 22432
rect 10597 22423 10655 22429
rect 10597 22420 10609 22423
rect 10468 22392 10609 22420
rect 10468 22380 10474 22392
rect 10597 22389 10609 22392
rect 10643 22389 10655 22423
rect 10597 22383 10655 22389
rect 10686 22380 10692 22432
rect 10744 22420 10750 22432
rect 11330 22420 11336 22432
rect 10744 22392 11336 22420
rect 10744 22380 10750 22392
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 11517 22423 11575 22429
rect 11517 22389 11529 22423
rect 11563 22420 11575 22423
rect 11882 22420 11888 22432
rect 11563 22392 11888 22420
rect 11563 22389 11575 22392
rect 11517 22383 11575 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 11977 22423 12035 22429
rect 11977 22389 11989 22423
rect 12023 22420 12035 22423
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 12023 22392 12173 22420
rect 12023 22389 12035 22392
rect 11977 22383 12035 22389
rect 12161 22389 12173 22392
rect 12207 22420 12219 22423
rect 12250 22420 12256 22432
rect 12207 22392 12256 22420
rect 12207 22389 12219 22392
rect 12161 22383 12219 22389
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 13262 22380 13268 22432
rect 13320 22420 13326 22432
rect 14642 22420 14648 22432
rect 13320 22392 14648 22420
rect 13320 22380 13326 22392
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 16758 22380 16764 22432
rect 16816 22380 16822 22432
rect 20625 22423 20683 22429
rect 20625 22389 20637 22423
rect 20671 22420 20683 22423
rect 20714 22420 20720 22432
rect 20671 22392 20720 22420
rect 20671 22389 20683 22392
rect 20625 22383 20683 22389
rect 20714 22380 20720 22392
rect 20772 22420 20778 22432
rect 21542 22420 21548 22432
rect 20772 22392 21548 22420
rect 20772 22380 20778 22392
rect 21542 22380 21548 22392
rect 21600 22380 21606 22432
rect 1104 22330 26864 22352
rect 1104 22278 4169 22330
rect 4221 22278 4233 22330
rect 4285 22278 4297 22330
rect 4349 22278 4361 22330
rect 4413 22278 4425 22330
rect 4477 22278 10608 22330
rect 10660 22278 10672 22330
rect 10724 22278 10736 22330
rect 10788 22278 10800 22330
rect 10852 22278 10864 22330
rect 10916 22278 17047 22330
rect 17099 22278 17111 22330
rect 17163 22278 17175 22330
rect 17227 22278 17239 22330
rect 17291 22278 17303 22330
rect 17355 22278 23486 22330
rect 23538 22278 23550 22330
rect 23602 22278 23614 22330
rect 23666 22278 23678 22330
rect 23730 22278 23742 22330
rect 23794 22278 26864 22330
rect 1104 22256 26864 22278
rect 4338 22176 4344 22228
rect 4396 22216 4402 22228
rect 4617 22219 4675 22225
rect 4617 22216 4629 22219
rect 4396 22188 4629 22216
rect 4396 22176 4402 22188
rect 4617 22185 4629 22188
rect 4663 22216 4675 22219
rect 4706 22216 4712 22228
rect 4663 22188 4712 22216
rect 4663 22185 4675 22188
rect 4617 22179 4675 22185
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 9122 22176 9128 22228
rect 9180 22176 9186 22228
rect 9585 22219 9643 22225
rect 9585 22185 9597 22219
rect 9631 22216 9643 22219
rect 9858 22216 9864 22228
rect 9631 22188 9864 22216
rect 9631 22185 9643 22188
rect 9585 22179 9643 22185
rect 9858 22176 9864 22188
rect 9916 22176 9922 22228
rect 9950 22176 9956 22228
rect 10008 22176 10014 22228
rect 10318 22176 10324 22228
rect 10376 22216 10382 22228
rect 10594 22216 10600 22228
rect 10376 22188 10600 22216
rect 10376 22176 10382 22188
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 11146 22176 11152 22228
rect 11204 22216 11210 22228
rect 11241 22219 11299 22225
rect 11241 22216 11253 22219
rect 11204 22188 11253 22216
rect 11204 22176 11210 22188
rect 11241 22185 11253 22188
rect 11287 22185 11299 22219
rect 11241 22179 11299 22185
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 12434 22216 12440 22228
rect 11388 22188 12440 22216
rect 11388 22176 11394 22188
rect 12434 22176 12440 22188
rect 12492 22176 12498 22228
rect 12526 22176 12532 22228
rect 12584 22216 12590 22228
rect 13262 22216 13268 22228
rect 12584 22188 13268 22216
rect 12584 22176 12590 22188
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 14182 22176 14188 22228
rect 14240 22176 14246 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 16758 22216 16764 22228
rect 16632 22188 16764 22216
rect 16632 22176 16638 22188
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 18506 22176 18512 22228
rect 18564 22176 18570 22228
rect 18966 22176 18972 22228
rect 19024 22176 19030 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 19245 22219 19303 22225
rect 19245 22216 19257 22219
rect 19116 22188 19257 22216
rect 19116 22176 19122 22188
rect 19245 22185 19257 22188
rect 19291 22185 19303 22219
rect 19245 22179 19303 22185
rect 19628 22188 19840 22216
rect 4172 22120 5120 22148
rect 3344 22052 4016 22080
rect 3344 22024 3372 22052
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 2866 22012 2872 22024
rect 2464 21984 2872 22012
rect 2464 21972 2470 21984
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 3145 22015 3203 22021
rect 3145 21981 3157 22015
rect 3191 21981 3203 22015
rect 3145 21975 3203 21981
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 21981 3295 22015
rect 3237 21975 3295 21981
rect 1578 21836 1584 21888
rect 1636 21836 1642 21888
rect 2498 21836 2504 21888
rect 2556 21836 2562 21888
rect 2774 21836 2780 21888
rect 2832 21836 2838 21888
rect 2958 21836 2964 21888
rect 3016 21836 3022 21888
rect 3160 21876 3188 21975
rect 3252 21944 3280 21975
rect 3326 21972 3332 22024
rect 3384 21972 3390 22024
rect 3988 22021 4016 22052
rect 4172 22024 4200 22120
rect 5092 22080 5120 22120
rect 9490 22108 9496 22160
rect 9548 22148 9554 22160
rect 9968 22148 9996 22176
rect 9548 22120 11560 22148
rect 9548 22108 9554 22120
rect 11532 22092 11560 22120
rect 11606 22108 11612 22160
rect 11664 22108 11670 22160
rect 12066 22148 12072 22160
rect 11808 22120 12072 22148
rect 6270 22080 6276 22092
rect 4264 22052 5028 22080
rect 5092 22052 5764 22080
rect 3421 22015 3479 22021
rect 3421 21981 3433 22015
rect 3467 22012 3479 22015
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 3467 21984 3801 22012
rect 3467 21981 3479 21984
rect 3421 21975 3479 21981
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4062 21972 4068 22024
rect 4120 21972 4126 22024
rect 4154 21972 4160 22024
rect 4212 21972 4218 22024
rect 4264 22021 4292 22052
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 21981 4307 22015
rect 4893 22015 4951 22021
rect 4893 22012 4905 22015
rect 4249 21975 4307 21981
rect 4448 21984 4905 22012
rect 3510 21944 3516 21956
rect 3252 21916 3516 21944
rect 3510 21904 3516 21916
rect 3568 21944 3574 21956
rect 4080 21944 4108 21972
rect 4448 21944 4476 21984
rect 3568 21916 4108 21944
rect 4264 21916 4476 21944
rect 4571 21981 4629 21984
rect 4571 21947 4583 21981
rect 4617 21947 4629 21981
rect 4893 21981 4905 21984
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 4571 21941 4629 21947
rect 4801 21947 4859 21953
rect 3568 21904 3574 21916
rect 3694 21876 3700 21888
rect 3160 21848 3700 21876
rect 3694 21836 3700 21848
rect 3752 21876 3758 21888
rect 4264 21876 4292 21916
rect 4801 21913 4813 21947
rect 4847 21944 4859 21947
rect 5000 21944 5028 22052
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5169 22015 5227 22021
rect 5169 22012 5181 22015
rect 5132 21984 5181 22012
rect 5132 21972 5138 21984
rect 5169 21981 5181 21984
rect 5215 21981 5227 22015
rect 5169 21975 5227 21981
rect 5534 21972 5540 22024
rect 5592 21972 5598 22024
rect 5736 22021 5764 22052
rect 5920 22052 6276 22080
rect 5920 22024 5948 22052
rect 6270 22040 6276 22052
rect 6328 22040 6334 22092
rect 9122 22040 9128 22092
rect 9180 22080 9186 22092
rect 9180 22052 9628 22080
rect 9180 22040 9186 22052
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 5442 21944 5448 21956
rect 4847 21916 5448 21944
rect 4847 21913 4859 21916
rect 4801 21907 4859 21913
rect 5442 21904 5448 21916
rect 5500 21904 5506 21956
rect 3752 21848 4292 21876
rect 3752 21836 3758 21848
rect 4430 21836 4436 21888
rect 4488 21836 4494 21888
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 4985 21879 5043 21885
rect 4985 21876 4997 21879
rect 4764 21848 4997 21876
rect 4764 21836 4770 21848
rect 4985 21845 4997 21848
rect 5031 21845 5043 21879
rect 4985 21839 5043 21845
rect 5258 21836 5264 21888
rect 5316 21836 5322 21888
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 5629 21879 5687 21885
rect 5629 21876 5641 21879
rect 5408 21848 5641 21876
rect 5408 21836 5414 21848
rect 5629 21845 5641 21848
rect 5675 21845 5687 21879
rect 5736 21876 5764 21975
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9398 22012 9404 22024
rect 8444 21984 9404 22012
rect 8444 21972 8450 21984
rect 6178 21904 6184 21956
rect 6236 21904 6242 21956
rect 7190 21904 7196 21956
rect 7248 21904 7254 21956
rect 8956 21953 8984 21984
rect 9398 21972 9404 21984
rect 9456 21972 9462 22024
rect 9600 22021 9628 22052
rect 11514 22040 11520 22092
rect 11572 22040 11578 22092
rect 11624 22080 11652 22108
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 11624 22052 11713 22080
rect 11701 22049 11713 22052
rect 11747 22049 11759 22083
rect 11701 22043 11759 22049
rect 9585 22015 9643 22021
rect 9585 21981 9597 22015
rect 9631 21981 9643 22015
rect 9585 21975 9643 21981
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 10008 21984 11437 22012
rect 10008 21972 10014 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11606 21972 11612 22024
rect 11664 22012 11670 22024
rect 11808 22012 11836 22120
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 18984 22148 19012 22176
rect 19628 22148 19656 22188
rect 18984 22120 19656 22148
rect 19812 22148 19840 22188
rect 20070 22176 20076 22228
rect 20128 22176 20134 22228
rect 20530 22176 20536 22228
rect 20588 22176 20594 22228
rect 21269 22219 21327 22225
rect 21269 22185 21281 22219
rect 21315 22216 21327 22219
rect 21358 22216 21364 22228
rect 21315 22188 21364 22216
rect 21315 22185 21327 22188
rect 21269 22179 21327 22185
rect 21358 22176 21364 22188
rect 21416 22176 21422 22228
rect 20088 22148 20116 22176
rect 21634 22148 21640 22160
rect 19812 22120 21640 22148
rect 16390 22080 16396 22092
rect 11664 21984 11836 22012
rect 11900 22052 16396 22080
rect 11664 21972 11670 21984
rect 8941 21947 8999 21953
rect 8941 21913 8953 21947
rect 8987 21944 8999 21947
rect 8987 21916 9021 21944
rect 8987 21913 8999 21916
rect 8941 21907 8999 21913
rect 9490 21904 9496 21956
rect 9548 21944 9554 21956
rect 9769 21947 9827 21953
rect 9769 21944 9781 21947
rect 9548 21916 9781 21944
rect 9548 21904 9554 21916
rect 9769 21913 9781 21916
rect 9815 21944 9827 21947
rect 9858 21944 9864 21956
rect 9815 21916 9864 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 10226 21944 10232 21956
rect 9968 21916 10232 21944
rect 6454 21876 6460 21888
rect 5736 21848 6460 21876
rect 5629 21839 5687 21845
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 6880 21848 7665 21876
rect 6880 21836 6886 21848
rect 7653 21845 7665 21848
rect 7699 21876 7711 21879
rect 9141 21879 9199 21885
rect 9141 21876 9153 21879
rect 7699 21848 9153 21876
rect 7699 21845 7711 21848
rect 7653 21839 7711 21845
rect 9141 21845 9153 21848
rect 9187 21845 9199 21879
rect 9141 21839 9199 21845
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9674 21876 9680 21888
rect 9355 21848 9680 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 9968 21885 9996 21916
rect 10226 21904 10232 21916
rect 10284 21904 10290 21956
rect 10502 21904 10508 21956
rect 10560 21944 10566 21956
rect 11900 21944 11928 22052
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 16485 22083 16543 22089
rect 16485 22049 16497 22083
rect 16531 22080 16543 22083
rect 16850 22080 16856 22092
rect 16531 22052 16856 22080
rect 16531 22049 16543 22052
rect 16485 22043 16543 22049
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 17221 22083 17279 22089
rect 17221 22049 17233 22083
rect 17267 22080 17279 22083
rect 17954 22080 17960 22092
rect 17267 22052 17960 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 19628 22089 19656 22120
rect 21634 22108 21640 22120
rect 21692 22108 21698 22160
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 18800 22052 19533 22080
rect 18800 22024 18828 22052
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 19521 22043 19579 22049
rect 19613 22083 19671 22089
rect 19613 22049 19625 22083
rect 19659 22049 19671 22083
rect 19613 22043 19671 22049
rect 19706 22083 19764 22089
rect 19706 22049 19718 22083
rect 19752 22080 19764 22083
rect 19886 22080 19892 22092
rect 19752 22052 19892 22080
rect 19752 22049 19764 22052
rect 19706 22043 19764 22049
rect 12250 21972 12256 22024
rect 12308 21972 12314 22024
rect 15930 21972 15936 22024
rect 15988 21972 15994 22024
rect 16577 22015 16635 22021
rect 16577 21981 16589 22015
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 10560 21916 11928 21944
rect 12069 21947 12127 21953
rect 10560 21904 10566 21916
rect 12069 21913 12081 21947
rect 12115 21944 12127 21947
rect 12115 21916 12434 21944
rect 12115 21913 12127 21916
rect 12069 21907 12127 21913
rect 9968 21879 10027 21885
rect 9968 21848 9981 21879
rect 9969 21845 9981 21848
rect 10015 21845 10027 21879
rect 9969 21839 10027 21845
rect 10134 21836 10140 21888
rect 10192 21836 10198 21888
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 11020 21848 11897 21876
rect 11020 21836 11026 21848
rect 11885 21845 11897 21848
rect 11931 21845 11943 21879
rect 12406 21876 12434 21916
rect 15194 21904 15200 21956
rect 15252 21904 15258 21956
rect 15654 21904 15660 21956
rect 15712 21904 15718 21956
rect 16592 21944 16620 21975
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 17129 22015 17187 22021
rect 17129 22012 17141 22015
rect 16816 21984 17141 22012
rect 16816 21972 16822 21984
rect 17129 21981 17141 21984
rect 17175 22012 17187 22015
rect 17586 22012 17592 22024
rect 17175 21984 17592 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 18104 21984 18153 22012
rect 18104 21972 18110 21984
rect 18141 21981 18153 21984
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 17497 21947 17555 21953
rect 17497 21944 17509 21947
rect 16592 21916 17509 21944
rect 17497 21913 17509 21916
rect 17543 21913 17555 21947
rect 18156 21944 18184 21975
rect 18690 21972 18696 22024
rect 18748 21972 18754 22024
rect 18782 21972 18788 22024
rect 18840 21972 18846 22024
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19536 22012 19564 22043
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20806 22080 20812 22092
rect 19996 22052 20812 22080
rect 19996 22012 20024 22052
rect 20806 22040 20812 22052
rect 20864 22080 20870 22092
rect 20901 22083 20959 22089
rect 20901 22080 20913 22083
rect 20864 22052 20913 22080
rect 20864 22040 20870 22052
rect 20901 22049 20913 22052
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 21542 22040 21548 22092
rect 21600 22040 21606 22092
rect 22646 22040 22652 22092
rect 22704 22040 22710 22092
rect 19536 21984 20024 22012
rect 19429 21975 19487 21981
rect 18598 21944 18604 21956
rect 18156 21916 18604 21944
rect 17497 21907 17555 21913
rect 18598 21904 18604 21916
rect 18656 21944 18662 21956
rect 18969 21947 19027 21953
rect 18969 21944 18981 21947
rect 18656 21916 18981 21944
rect 18656 21904 18662 21916
rect 18969 21913 18981 21916
rect 19015 21944 19027 21947
rect 19444 21944 19472 21975
rect 20070 21972 20076 22024
rect 20128 21972 20134 22024
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20717 22015 20775 22021
rect 20717 22012 20729 22015
rect 20680 21984 20729 22012
rect 20680 21972 20686 21984
rect 20717 21981 20729 21984
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 21634 21972 21640 22024
rect 21692 21972 21698 22024
rect 22554 21972 22560 22024
rect 22612 21972 22618 22024
rect 20640 21944 20668 21972
rect 22572 21944 22600 21972
rect 19015 21916 20668 21944
rect 22066 21916 22600 21944
rect 19015 21913 19027 21916
rect 18969 21907 19027 21913
rect 18230 21876 18236 21888
rect 12406 21848 18236 21876
rect 11885 21839 11943 21845
rect 18230 21836 18236 21848
rect 18288 21876 18294 21888
rect 18690 21876 18696 21888
rect 18288 21848 18696 21876
rect 18288 21836 18294 21848
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19978 21836 19984 21888
rect 20036 21836 20042 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 22066 21876 22094 21916
rect 20128 21848 22094 21876
rect 20128 21836 20134 21848
rect 1104 21786 26864 21808
rect 1104 21734 4829 21786
rect 4881 21734 4893 21786
rect 4945 21734 4957 21786
rect 5009 21734 5021 21786
rect 5073 21734 5085 21786
rect 5137 21734 11268 21786
rect 11320 21734 11332 21786
rect 11384 21734 11396 21786
rect 11448 21734 11460 21786
rect 11512 21734 11524 21786
rect 11576 21734 17707 21786
rect 17759 21734 17771 21786
rect 17823 21734 17835 21786
rect 17887 21734 17899 21786
rect 17951 21734 17963 21786
rect 18015 21734 24146 21786
rect 24198 21734 24210 21786
rect 24262 21734 24274 21786
rect 24326 21734 24338 21786
rect 24390 21734 24402 21786
rect 24454 21734 26864 21786
rect 1104 21712 26864 21734
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 3786 21672 3792 21684
rect 3384 21644 3792 21672
rect 3384 21632 3390 21644
rect 3436 21613 3464 21644
rect 3786 21632 3792 21644
rect 3844 21632 3850 21684
rect 4249 21675 4307 21681
rect 4249 21672 4261 21675
rect 3896 21644 4261 21672
rect 3421 21607 3479 21613
rect 3421 21573 3433 21607
rect 3467 21573 3479 21607
rect 3421 21567 3479 21573
rect 3510 21564 3516 21616
rect 3568 21604 3574 21616
rect 3896 21613 3924 21644
rect 4249 21641 4261 21644
rect 4295 21641 4307 21675
rect 4249 21635 4307 21641
rect 5537 21675 5595 21681
rect 5537 21641 5549 21675
rect 5583 21672 5595 21675
rect 6178 21672 6184 21684
rect 5583 21644 6184 21672
rect 5583 21641 5595 21644
rect 5537 21635 5595 21641
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 6454 21632 6460 21684
rect 6512 21632 6518 21684
rect 7101 21675 7159 21681
rect 7101 21641 7113 21675
rect 7147 21672 7159 21675
rect 7190 21672 7196 21684
rect 7147 21644 7196 21672
rect 7147 21641 7159 21644
rect 7101 21635 7159 21641
rect 7190 21632 7196 21644
rect 7248 21632 7254 21684
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 10226 21672 10232 21684
rect 8260 21644 10232 21672
rect 8260 21632 8266 21644
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 14642 21632 14648 21684
rect 14700 21632 14706 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 15289 21675 15347 21681
rect 15289 21672 15301 21675
rect 15252 21644 15301 21672
rect 15252 21632 15258 21644
rect 15289 21641 15301 21644
rect 15335 21641 15347 21675
rect 15289 21635 15347 21641
rect 15654 21632 15660 21684
rect 15712 21632 15718 21684
rect 18233 21675 18291 21681
rect 18233 21641 18245 21675
rect 18279 21672 18291 21675
rect 18322 21672 18328 21684
rect 18279 21644 18328 21672
rect 18279 21641 18291 21644
rect 18233 21635 18291 21641
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 3881 21607 3939 21613
rect 3568 21576 3832 21604
rect 3568 21564 3574 21576
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 3804 21545 3832 21576
rect 3881 21573 3893 21607
rect 3927 21573 3939 21607
rect 4706 21604 4712 21616
rect 3881 21567 3939 21573
rect 4540 21576 4712 21604
rect 3671 21539 3729 21545
rect 3671 21505 3683 21539
rect 3717 21536 3729 21539
rect 3789 21539 3847 21545
rect 3717 21505 3740 21536
rect 3671 21499 3740 21505
rect 3789 21505 3801 21539
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 1719 21440 2774 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 2746 21400 2774 21440
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 3712 21468 3740 21499
rect 3970 21496 3976 21548
rect 4028 21496 4034 21548
rect 4540 21545 4568 21576
rect 4706 21564 4712 21576
rect 4764 21564 4770 21616
rect 6917 21607 6975 21613
rect 6917 21604 6929 21607
rect 5644 21576 6929 21604
rect 4525 21539 4583 21545
rect 4525 21505 4537 21539
rect 4571 21505 4583 21539
rect 4801 21539 4859 21545
rect 4801 21536 4813 21539
rect 4525 21499 4583 21505
rect 4632 21508 4813 21536
rect 3878 21468 3884 21480
rect 3712 21440 3884 21468
rect 3878 21428 3884 21440
rect 3936 21468 3942 21480
rect 3936 21440 4292 21468
rect 3936 21428 3942 21440
rect 4157 21403 4215 21409
rect 4157 21400 4169 21403
rect 2746 21372 4169 21400
rect 4157 21369 4169 21372
rect 4203 21369 4215 21403
rect 4264 21400 4292 21440
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 4632 21468 4660 21508
rect 4801 21505 4813 21508
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21505 5043 21539
rect 5169 21539 5227 21545
rect 5169 21538 5181 21539
rect 5215 21538 5227 21539
rect 5261 21539 5319 21545
rect 4985 21499 5043 21505
rect 4396 21440 4660 21468
rect 4396 21428 4402 21440
rect 4706 21428 4712 21480
rect 4764 21468 4770 21480
rect 5000 21468 5028 21499
rect 5166 21486 5172 21538
rect 5224 21486 5230 21538
rect 5261 21505 5273 21539
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 4764 21440 5028 21468
rect 4764 21428 4770 21440
rect 5276 21400 5304 21499
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 5644 21468 5672 21576
rect 6917 21573 6929 21576
rect 6963 21604 6975 21607
rect 8220 21604 8248 21632
rect 6963 21576 8248 21604
rect 12253 21607 12311 21613
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 12253 21573 12265 21607
rect 12299 21604 12311 21607
rect 12434 21604 12440 21616
rect 12299 21576 12440 21604
rect 12299 21573 12311 21576
rect 12253 21567 12311 21573
rect 12434 21564 12440 21576
rect 12492 21564 12498 21616
rect 13538 21564 13544 21616
rect 13596 21564 13602 21616
rect 15930 21604 15936 21616
rect 14292 21576 15936 21604
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 6089 21539 6147 21545
rect 6089 21536 6101 21539
rect 5776 21508 6101 21536
rect 5776 21496 5782 21508
rect 6089 21505 6101 21508
rect 6135 21536 6147 21539
rect 6641 21539 6699 21545
rect 6641 21536 6653 21539
rect 6135 21508 6653 21536
rect 6135 21505 6147 21508
rect 6089 21499 6147 21505
rect 6641 21505 6653 21508
rect 6687 21536 6699 21539
rect 6822 21536 6828 21548
rect 6687 21508 6828 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 7098 21496 7104 21548
rect 7156 21536 7162 21548
rect 14292 21545 14320 21576
rect 15930 21564 15936 21576
rect 15988 21604 15994 21616
rect 16758 21604 16764 21616
rect 15988 21576 16764 21604
rect 15988 21564 15994 21576
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 18966 21604 18972 21616
rect 17788 21576 18972 21604
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 7156 21508 7205 21536
rect 7156 21496 7162 21508
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 14458 21496 14464 21548
rect 14516 21536 14522 21548
rect 14737 21539 14795 21545
rect 14737 21536 14749 21539
rect 14516 21508 14749 21536
rect 14516 21496 14522 21508
rect 14737 21505 14749 21508
rect 14783 21505 14795 21539
rect 14737 21499 14795 21505
rect 15286 21496 15292 21548
rect 15344 21536 15350 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 15344 21508 15393 21536
rect 15344 21496 15350 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 5813 21471 5871 21477
rect 5813 21468 5825 21471
rect 5644 21440 5825 21468
rect 5813 21437 5825 21440
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21437 5963 21471
rect 5905 21431 5963 21437
rect 5920 21400 5948 21431
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 6546 21468 6552 21480
rect 6052 21440 6552 21468
rect 6052 21428 6058 21440
rect 6546 21428 6552 21440
rect 6604 21428 6610 21480
rect 6733 21471 6791 21477
rect 6733 21468 6745 21471
rect 6656 21440 6745 21468
rect 6454 21400 6460 21412
rect 4264 21372 5304 21400
rect 5828 21372 6460 21400
rect 4157 21363 4215 21369
rect 5828 21344 5856 21372
rect 6454 21360 6460 21372
rect 6512 21400 6518 21412
rect 6656 21400 6684 21440
rect 6733 21437 6745 21440
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 13998 21428 14004 21480
rect 14056 21428 14062 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 15488 21468 15516 21499
rect 16390 21496 16396 21548
rect 16448 21536 16454 21548
rect 17788 21545 17816 21576
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 16448 21508 17785 21536
rect 16448 21496 16454 21508
rect 17773 21505 17785 21508
rect 17819 21505 17831 21539
rect 17773 21499 17831 21505
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 15120 21440 15516 21468
rect 15120 21409 15148 21440
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 20070 21468 20076 21480
rect 17644 21440 20076 21468
rect 17644 21428 17650 21440
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 6512 21372 6684 21400
rect 15105 21403 15163 21409
rect 6512 21360 6518 21372
rect 15105 21369 15117 21403
rect 15151 21369 15163 21403
rect 15105 21363 15163 21369
rect 3786 21292 3792 21344
rect 3844 21332 3850 21344
rect 4338 21332 4344 21344
rect 3844 21304 4344 21332
rect 3844 21292 3850 21304
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 4709 21335 4767 21341
rect 4709 21301 4721 21335
rect 4755 21332 4767 21335
rect 4890 21332 4896 21344
rect 4755 21304 4896 21332
rect 4755 21301 4767 21304
rect 4709 21295 4767 21301
rect 4890 21292 4896 21304
rect 4948 21332 4954 21344
rect 5350 21332 5356 21344
rect 4948 21304 5356 21332
rect 4948 21292 4954 21304
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 5626 21292 5632 21344
rect 5684 21292 5690 21344
rect 5810 21292 5816 21344
rect 5868 21292 5874 21344
rect 6822 21292 6828 21344
rect 6880 21292 6886 21344
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 17911 21335 17969 21341
rect 17911 21332 17923 21335
rect 13320 21304 17923 21332
rect 13320 21292 13326 21304
rect 17911 21301 17923 21304
rect 17957 21332 17969 21335
rect 18782 21332 18788 21344
rect 17957 21304 18788 21332
rect 17957 21301 17969 21304
rect 17911 21295 17969 21301
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 1104 21242 26864 21264
rect 1104 21190 4169 21242
rect 4221 21190 4233 21242
rect 4285 21190 4297 21242
rect 4349 21190 4361 21242
rect 4413 21190 4425 21242
rect 4477 21190 10608 21242
rect 10660 21190 10672 21242
rect 10724 21190 10736 21242
rect 10788 21190 10800 21242
rect 10852 21190 10864 21242
rect 10916 21190 17047 21242
rect 17099 21190 17111 21242
rect 17163 21190 17175 21242
rect 17227 21190 17239 21242
rect 17291 21190 17303 21242
rect 17355 21190 23486 21242
rect 23538 21190 23550 21242
rect 23602 21190 23614 21242
rect 23666 21190 23678 21242
rect 23730 21190 23742 21242
rect 23794 21190 26864 21242
rect 1104 21168 26864 21190
rect 3878 21088 3884 21140
rect 3936 21088 3942 21140
rect 4890 21128 4896 21140
rect 4080 21100 4896 21128
rect 3375 21063 3433 21069
rect 3375 21029 3387 21063
rect 3421 21060 3433 21063
rect 4080 21060 4108 21100
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 5166 21088 5172 21140
rect 5224 21088 5230 21140
rect 5350 21088 5356 21140
rect 5408 21128 5414 21140
rect 9950 21128 9956 21140
rect 5408 21100 9956 21128
rect 5408 21088 5414 21100
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 13081 21131 13139 21137
rect 13081 21097 13093 21131
rect 13127 21128 13139 21131
rect 13998 21128 14004 21140
rect 13127 21100 14004 21128
rect 13127 21097 13139 21100
rect 13081 21091 13139 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 16942 21088 16948 21140
rect 17000 21088 17006 21140
rect 3421 21032 4108 21060
rect 3421 21029 3433 21032
rect 3375 21023 3433 21029
rect 1394 20952 1400 21004
rect 1452 20992 1458 21004
rect 1581 20995 1639 21001
rect 1581 20992 1593 20995
rect 1452 20964 1593 20992
rect 1452 20952 1458 20964
rect 1581 20961 1593 20964
rect 1627 20961 1639 20995
rect 1581 20955 1639 20961
rect 1949 20995 2007 21001
rect 1949 20961 1961 20995
rect 1995 20992 2007 20995
rect 2958 20992 2964 21004
rect 1995 20964 2964 20992
rect 1995 20961 2007 20964
rect 1949 20955 2007 20961
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 4080 20933 4108 21032
rect 4154 21020 4160 21072
rect 4212 21060 4218 21072
rect 4249 21063 4307 21069
rect 4249 21060 4261 21063
rect 4212 21032 4261 21060
rect 4212 21020 4218 21032
rect 4249 21029 4261 21032
rect 4295 21029 4307 21063
rect 5258 21060 5264 21072
rect 4249 21023 4307 21029
rect 4632 21032 5264 21060
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 4341 20927 4399 20933
rect 4341 20893 4353 20927
rect 4387 20924 4399 20927
rect 4632 20924 4660 21032
rect 5258 21020 5264 21032
rect 5316 21020 5322 21072
rect 10318 21020 10324 21072
rect 10376 21020 10382 21072
rect 13538 21020 13544 21072
rect 13596 21060 13602 21072
rect 13817 21063 13875 21069
rect 13817 21060 13829 21063
rect 13596 21032 13829 21060
rect 13596 21020 13602 21032
rect 13817 21029 13829 21032
rect 13863 21029 13875 21063
rect 13817 21023 13875 21029
rect 5626 20992 5632 21004
rect 4724 20964 5632 20992
rect 4724 20933 4752 20964
rect 5626 20952 5632 20964
rect 5684 20952 5690 21004
rect 8938 20952 8944 21004
rect 8996 20952 9002 21004
rect 9125 20995 9183 21001
rect 9125 20961 9137 20995
rect 9171 20992 9183 20995
rect 9398 20992 9404 21004
rect 9171 20964 9404 20992
rect 9171 20961 9183 20964
rect 9125 20955 9183 20961
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 10336 20992 10364 21020
rect 10152 20964 10364 20992
rect 4387 20896 4660 20924
rect 4709 20927 4767 20933
rect 4387 20893 4399 20896
rect 4341 20887 4399 20893
rect 4709 20893 4721 20927
rect 4755 20893 4767 20927
rect 4709 20887 4767 20893
rect 2498 20816 2504 20868
rect 2556 20816 2562 20868
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 4172 20856 4200 20887
rect 4798 20884 4804 20936
rect 4856 20884 4862 20936
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20924 5043 20927
rect 5350 20924 5356 20936
rect 5031 20896 5356 20924
rect 5031 20893 5043 20896
rect 4985 20887 5043 20893
rect 3844 20828 4200 20856
rect 3844 20816 3850 20828
rect 4614 20816 4620 20868
rect 4672 20856 4678 20868
rect 5000 20856 5028 20887
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 9217 20927 9275 20933
rect 9217 20893 9229 20927
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 4672 20828 5028 20856
rect 4672 20816 4678 20828
rect 7006 20816 7012 20868
rect 7064 20816 7070 20868
rect 9030 20816 9036 20868
rect 9088 20856 9094 20868
rect 9232 20856 9260 20887
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 10152 20933 10180 20964
rect 13446 20952 13452 21004
rect 13504 20992 13510 21004
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 13504 20964 14565 20992
rect 13504 20952 13510 20964
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 10137 20927 10195 20933
rect 10137 20924 10149 20927
rect 9732 20896 10149 20924
rect 9732 20884 9738 20896
rect 10137 20893 10149 20896
rect 10183 20893 10195 20927
rect 10137 20887 10195 20893
rect 10226 20884 10232 20936
rect 10284 20884 10290 20936
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 10376 20896 10425 20924
rect 10376 20884 10382 20896
rect 10413 20893 10425 20896
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 13909 20927 13967 20933
rect 13909 20893 13921 20927
rect 13955 20924 13967 20927
rect 15286 20924 15292 20936
rect 13955 20896 15292 20924
rect 13955 20893 13967 20896
rect 13909 20887 13967 20893
rect 9088 20828 9260 20856
rect 9088 20816 9094 20828
rect 9950 20816 9956 20868
rect 10008 20816 10014 20868
rect 12912 20856 12940 20887
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 12912 20828 14136 20856
rect 5721 20791 5779 20797
rect 5721 20757 5733 20791
rect 5767 20788 5779 20791
rect 5902 20788 5908 20800
rect 5767 20760 5908 20788
rect 5767 20757 5779 20760
rect 5721 20751 5779 20757
rect 5902 20748 5908 20760
rect 5960 20788 5966 20800
rect 6454 20788 6460 20800
rect 5960 20760 6460 20788
rect 5960 20748 5966 20760
rect 6454 20748 6460 20760
rect 6512 20748 6518 20800
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 8941 20791 8999 20797
rect 8941 20788 8953 20791
rect 8720 20760 8953 20788
rect 8720 20748 8726 20760
rect 8941 20757 8953 20760
rect 8987 20757 8999 20791
rect 8941 20751 8999 20757
rect 9766 20748 9772 20800
rect 9824 20748 9830 20800
rect 9858 20748 9864 20800
rect 9916 20788 9922 20800
rect 14108 20797 14136 20828
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 15102 20856 15108 20868
rect 14516 20828 15108 20856
rect 14516 20816 14522 20828
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 15654 20816 15660 20868
rect 15712 20816 15718 20868
rect 10229 20791 10287 20797
rect 10229 20788 10241 20791
rect 9916 20760 10241 20788
rect 9916 20748 9922 20760
rect 10229 20757 10241 20760
rect 10275 20757 10287 20791
rect 10229 20751 10287 20757
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 17589 20791 17647 20797
rect 17589 20788 17601 20791
rect 17460 20760 17601 20788
rect 17460 20748 17466 20760
rect 17589 20757 17601 20760
rect 17635 20757 17647 20791
rect 17589 20751 17647 20757
rect 1104 20698 26864 20720
rect 1104 20646 4829 20698
rect 4881 20646 4893 20698
rect 4945 20646 4957 20698
rect 5009 20646 5021 20698
rect 5073 20646 5085 20698
rect 5137 20646 11268 20698
rect 11320 20646 11332 20698
rect 11384 20646 11396 20698
rect 11448 20646 11460 20698
rect 11512 20646 11524 20698
rect 11576 20646 17707 20698
rect 17759 20646 17771 20698
rect 17823 20646 17835 20698
rect 17887 20646 17899 20698
rect 17951 20646 17963 20698
rect 18015 20646 24146 20698
rect 24198 20646 24210 20698
rect 24262 20646 24274 20698
rect 24326 20646 24338 20698
rect 24390 20646 24402 20698
rect 24454 20646 26864 20698
rect 1104 20624 26864 20646
rect 3421 20587 3479 20593
rect 3421 20553 3433 20587
rect 3467 20584 3479 20587
rect 3510 20584 3516 20596
rect 3467 20556 3516 20584
rect 3467 20553 3479 20556
rect 3421 20547 3479 20553
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 4065 20587 4123 20593
rect 4065 20584 4077 20587
rect 4028 20556 4077 20584
rect 4028 20544 4034 20556
rect 4065 20553 4077 20556
rect 4111 20553 4123 20587
rect 4065 20547 4123 20553
rect 4706 20544 4712 20596
rect 4764 20584 4770 20596
rect 4893 20587 4951 20593
rect 4893 20584 4905 20587
rect 4764 20556 4905 20584
rect 4764 20544 4770 20556
rect 4893 20553 4905 20556
rect 4939 20553 4951 20587
rect 4893 20547 4951 20553
rect 5534 20544 5540 20596
rect 5592 20544 5598 20596
rect 8202 20584 8208 20596
rect 6380 20556 8208 20584
rect 3786 20516 3792 20528
rect 3068 20488 3792 20516
rect 3068 20457 3096 20488
rect 3786 20476 3792 20488
rect 3844 20516 3850 20528
rect 5166 20525 5172 20528
rect 3881 20519 3939 20525
rect 3881 20516 3893 20519
rect 3844 20488 3893 20516
rect 3844 20476 3850 20488
rect 3881 20485 3893 20488
rect 3927 20485 3939 20519
rect 3881 20479 3939 20485
rect 5153 20519 5172 20525
rect 5153 20485 5165 20519
rect 5153 20479 5172 20485
rect 5166 20476 5172 20479
rect 5224 20476 5230 20528
rect 5353 20519 5411 20525
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5399 20488 5488 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 3694 20408 3700 20460
rect 3752 20448 3758 20460
rect 5460 20457 5488 20488
rect 5626 20476 5632 20528
rect 5684 20516 5690 20528
rect 5684 20488 5948 20516
rect 5684 20476 5690 20488
rect 5445 20451 5503 20457
rect 3752 20420 4384 20448
rect 3752 20408 3758 20420
rect 3145 20383 3203 20389
rect 3145 20349 3157 20383
rect 3191 20380 3203 20383
rect 4154 20380 4160 20392
rect 3191 20352 4160 20380
rect 3191 20349 3203 20352
rect 3145 20343 3203 20349
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 3602 20272 3608 20324
rect 3660 20312 3666 20324
rect 4062 20312 4068 20324
rect 3660 20284 4068 20312
rect 3660 20272 3666 20284
rect 4062 20272 4068 20284
rect 4120 20312 4126 20324
rect 4264 20312 4292 20343
rect 4120 20284 4292 20312
rect 4356 20312 4384 20420
rect 5445 20417 5457 20451
rect 5491 20448 5503 20451
rect 5718 20448 5724 20460
rect 5491 20420 5724 20448
rect 5491 20417 5503 20420
rect 5445 20411 5503 20417
rect 5718 20408 5724 20420
rect 5776 20408 5782 20460
rect 5920 20457 5948 20488
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20448 5963 20451
rect 5994 20448 6000 20460
rect 5951 20420 6000 20448
rect 5951 20417 5963 20420
rect 5905 20411 5963 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20380 5687 20383
rect 6380 20380 6408 20556
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 9125 20587 9183 20593
rect 9125 20584 9137 20587
rect 8996 20556 9137 20584
rect 8996 20544 9002 20556
rect 9125 20553 9137 20556
rect 9171 20553 9183 20587
rect 9125 20547 9183 20553
rect 9309 20587 9367 20593
rect 9309 20553 9321 20587
rect 9355 20584 9367 20587
rect 9766 20584 9772 20596
rect 9355 20556 9772 20584
rect 9355 20553 9367 20556
rect 9309 20547 9367 20553
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10100 20556 10885 20584
rect 10100 20544 10106 20556
rect 7282 20476 7288 20528
rect 7340 20476 7346 20528
rect 6454 20408 6460 20460
rect 6512 20408 6518 20460
rect 8220 20448 8248 20544
rect 10152 20525 10180 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 11698 20584 11704 20596
rect 10873 20547 10931 20553
rect 11532 20556 11704 20584
rect 10137 20519 10195 20525
rect 10137 20485 10149 20519
rect 10183 20485 10195 20519
rect 10137 20479 10195 20485
rect 10244 20488 11008 20516
rect 8941 20451 8999 20457
rect 8941 20448 8953 20451
rect 8220 20420 8953 20448
rect 8941 20417 8953 20420
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 9950 20457 9956 20460
rect 9927 20451 9956 20457
rect 9732 20420 9812 20448
rect 9732 20408 9738 20420
rect 5675 20352 6408 20380
rect 5675 20349 5687 20352
rect 5629 20343 5687 20349
rect 4985 20315 5043 20321
rect 4985 20312 4997 20315
rect 4356 20284 4997 20312
rect 4120 20272 4126 20284
rect 4985 20281 4997 20284
rect 5031 20281 5043 20315
rect 4985 20275 5043 20281
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 5644 20312 5672 20343
rect 6730 20340 6736 20392
rect 6788 20340 6794 20392
rect 9784 20389 9812 20420
rect 9927 20417 9939 20451
rect 9927 20411 9956 20417
rect 9950 20408 9956 20411
rect 10008 20408 10014 20460
rect 10244 20457 10272 20488
rect 10980 20460 11008 20488
rect 11330 20476 11336 20528
rect 11388 20516 11394 20528
rect 11532 20525 11560 20556
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 17034 20544 17040 20596
rect 17092 20584 17098 20596
rect 24578 20584 24584 20596
rect 17092 20556 24584 20584
rect 17092 20544 17098 20556
rect 24578 20544 24584 20556
rect 24636 20544 24642 20596
rect 11517 20519 11575 20525
rect 11517 20516 11529 20519
rect 11388 20488 11529 20516
rect 11388 20476 11394 20488
rect 11517 20485 11529 20488
rect 11563 20485 11575 20519
rect 17402 20516 17408 20528
rect 11517 20479 11575 20485
rect 15488 20488 17408 20516
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10229 20451 10287 20457
rect 10091 20420 10180 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20349 9827 20383
rect 10152 20380 10180 20420
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10229 20411 10287 20417
rect 10336 20420 10701 20448
rect 10336 20380 10364 20420
rect 10689 20417 10701 20420
rect 10735 20448 10747 20451
rect 10870 20448 10876 20460
rect 10735 20420 10876 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 11790 20448 11796 20460
rect 11747 20420 11796 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 15488 20457 15516 20488
rect 17402 20476 17408 20488
rect 17460 20476 17466 20528
rect 18598 20516 18604 20528
rect 18446 20488 18604 20516
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18782 20476 18788 20528
rect 18840 20516 18846 20528
rect 18840 20488 19932 20516
rect 18840 20476 18846 20488
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 10152 20352 10364 20380
rect 9769 20343 9827 20349
rect 10502 20340 10508 20392
rect 10560 20380 10566 20392
rect 10560 20352 12434 20380
rect 10560 20340 10566 20352
rect 5500 20284 5672 20312
rect 9677 20315 9735 20321
rect 5500 20272 5506 20284
rect 9677 20281 9689 20315
rect 9723 20312 9735 20315
rect 10226 20312 10232 20324
rect 9723 20284 10232 20312
rect 9723 20281 9735 20284
rect 9677 20275 9735 20281
rect 10226 20272 10232 20284
rect 10284 20312 10290 20324
rect 10413 20315 10471 20321
rect 10413 20312 10425 20315
rect 10284 20284 10425 20312
rect 10284 20272 10290 20284
rect 10413 20281 10425 20284
rect 10459 20281 10471 20315
rect 12406 20312 12434 20352
rect 15378 20340 15384 20392
rect 15436 20340 15442 20392
rect 15580 20380 15608 20411
rect 15930 20408 15936 20460
rect 15988 20408 15994 20460
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16908 20420 16957 20448
rect 16908 20408 16914 20420
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 19904 20457 19932 20488
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 19889 20451 19947 20457
rect 17359 20420 17724 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 16482 20380 16488 20392
rect 15580 20352 16488 20380
rect 16482 20340 16488 20352
rect 16540 20340 16546 20392
rect 14458 20312 14464 20324
rect 12406 20284 14464 20312
rect 10413 20275 10471 20281
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 16390 20272 16396 20324
rect 16448 20272 16454 20324
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17144 20312 17172 20411
rect 17696 20392 17724 20420
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20380 17463 20383
rect 17494 20380 17500 20392
rect 17451 20352 17500 20380
rect 17451 20349 17463 20352
rect 17405 20343 17463 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 17678 20340 17684 20392
rect 17736 20340 17742 20392
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18877 20383 18935 20389
rect 18877 20380 18889 20383
rect 18472 20352 18889 20380
rect 18472 20340 18478 20352
rect 18877 20349 18889 20352
rect 18923 20349 18935 20383
rect 18877 20343 18935 20349
rect 19150 20340 19156 20392
rect 19208 20340 19214 20392
rect 17000 20284 17172 20312
rect 17000 20272 17006 20284
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 5169 20247 5227 20253
rect 5169 20244 5181 20247
rect 4580 20216 5181 20244
rect 4580 20204 4586 20216
rect 5169 20213 5181 20216
rect 5215 20244 5227 20247
rect 5626 20244 5632 20256
rect 5215 20216 5632 20244
rect 5215 20213 5227 20216
rect 5169 20207 5227 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 5810 20253 5816 20256
rect 5767 20247 5816 20253
rect 5767 20213 5779 20247
rect 5813 20213 5816 20247
rect 5767 20207 5816 20213
rect 5810 20204 5816 20207
rect 5868 20204 5874 20256
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 10318 20244 10324 20256
rect 9355 20216 10324 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 10318 20204 10324 20216
rect 10376 20244 10382 20256
rect 10505 20247 10563 20253
rect 10505 20244 10517 20247
rect 10376 20216 10517 20244
rect 10376 20204 10382 20216
rect 10505 20213 10517 20216
rect 10551 20213 10563 20247
rect 10505 20207 10563 20213
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11204 20216 11897 20244
rect 11204 20204 11210 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16172 20216 16681 20244
rect 16172 20204 16178 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 1104 20154 26864 20176
rect 1104 20102 4169 20154
rect 4221 20102 4233 20154
rect 4285 20102 4297 20154
rect 4349 20102 4361 20154
rect 4413 20102 4425 20154
rect 4477 20102 10608 20154
rect 10660 20102 10672 20154
rect 10724 20102 10736 20154
rect 10788 20102 10800 20154
rect 10852 20102 10864 20154
rect 10916 20102 17047 20154
rect 17099 20102 17111 20154
rect 17163 20102 17175 20154
rect 17227 20102 17239 20154
rect 17291 20102 17303 20154
rect 17355 20102 23486 20154
rect 23538 20102 23550 20154
rect 23602 20102 23614 20154
rect 23666 20102 23678 20154
rect 23730 20102 23742 20154
rect 23794 20102 26864 20154
rect 1104 20080 26864 20102
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6788 20012 6929 20040
rect 6788 20000 6794 20012
rect 6917 20009 6929 20012
rect 6963 20009 6975 20043
rect 6917 20003 6975 20009
rect 7282 20000 7288 20052
rect 7340 20000 7346 20052
rect 9398 20000 9404 20052
rect 9456 20000 9462 20052
rect 9582 20000 9588 20052
rect 9640 20040 9646 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 9640 20012 10977 20040
rect 9640 20000 9646 20012
rect 10965 20009 10977 20012
rect 11011 20009 11023 20043
rect 10965 20003 11023 20009
rect 9858 19972 9864 19984
rect 8772 19944 9864 19972
rect 8386 19904 8392 19916
rect 7024 19876 8392 19904
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4672 19808 4997 19836
rect 4672 19796 4678 19808
rect 4985 19805 4997 19808
rect 5031 19836 5043 19839
rect 5166 19836 5172 19848
rect 5031 19808 5172 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19836 5411 19839
rect 5442 19836 5448 19848
rect 5399 19808 5448 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 5810 19836 5816 19848
rect 5592 19808 5816 19836
rect 5592 19796 5598 19808
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 7024 19845 7052 19876
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 7156 19808 7205 19836
rect 7156 19796 7162 19808
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 8481 19799 8539 19805
rect 4706 19728 4712 19780
rect 4764 19768 4770 19780
rect 4801 19771 4859 19777
rect 4801 19768 4813 19771
rect 4764 19740 4813 19768
rect 4764 19728 4770 19740
rect 4801 19737 4813 19740
rect 4847 19737 4859 19771
rect 8496 19768 8524 19799
rect 8662 19796 8668 19848
rect 8720 19796 8726 19848
rect 8772 19845 8800 19944
rect 9858 19932 9864 19944
rect 9916 19932 9922 19984
rect 10980 19972 11008 20003
rect 11790 20000 11796 20052
rect 11848 20000 11854 20052
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20009 12219 20043
rect 12161 20003 12219 20009
rect 10980 19944 11744 19972
rect 10781 19907 10839 19913
rect 8864 19876 10088 19904
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19805 8815 19839
rect 8757 19799 8815 19805
rect 8864 19768 8892 19876
rect 9030 19796 9036 19848
rect 9088 19796 9094 19848
rect 10060 19845 10088 19876
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 11146 19904 11152 19916
rect 10827 19876 11152 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 11606 19904 11612 19916
rect 11440 19876 11612 19904
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 10045 19839 10103 19845
rect 9815 19808 9996 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 8496 19740 8892 19768
rect 4801 19731 4859 19737
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 8996 19740 9413 19768
rect 8996 19728 9002 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 9490 19728 9496 19780
rect 9548 19768 9554 19780
rect 9861 19771 9919 19777
rect 9861 19768 9873 19771
rect 9548 19740 9873 19768
rect 9548 19728 9554 19740
rect 9861 19737 9873 19740
rect 9907 19737 9919 19771
rect 9861 19731 9919 19737
rect 1578 19660 1584 19712
rect 1636 19660 1642 19712
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 4617 19703 4675 19709
rect 4617 19700 4629 19703
rect 3568 19672 4629 19700
rect 3568 19660 3574 19672
rect 4617 19669 4629 19672
rect 4663 19669 4675 19703
rect 4617 19663 4675 19669
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 8754 19700 8760 19712
rect 8343 19672 8760 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 9968 19700 9996 19808
rect 10045 19805 10057 19839
rect 10091 19805 10103 19839
rect 10045 19799 10103 19805
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 10410 19836 10416 19848
rect 10367 19808 10416 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 10060 19768 10088 19799
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 10870 19836 10876 19848
rect 10643 19808 10876 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 10060 19740 10793 19768
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 11072 19768 11100 19799
rect 11330 19796 11336 19848
rect 11388 19796 11394 19848
rect 11440 19845 11468 19876
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 11716 19845 11744 19944
rect 11425 19839 11483 19845
rect 11425 19805 11437 19839
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 11072 19740 11529 19768
rect 10781 19731 10839 19737
rect 11517 19737 11529 19740
rect 11563 19768 11575 19771
rect 11606 19768 11612 19780
rect 11563 19740 11612 19768
rect 11563 19737 11575 19740
rect 11517 19731 11575 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 12176 19768 12204 20003
rect 16114 20000 16120 20052
rect 16172 20000 16178 20052
rect 16482 20000 16488 20052
rect 16540 20000 16546 20052
rect 17678 20040 17684 20052
rect 16868 20012 17684 20040
rect 14829 19975 14887 19981
rect 14829 19941 14841 19975
rect 14875 19972 14887 19975
rect 16025 19975 16083 19981
rect 16025 19972 16037 19975
rect 14875 19944 16037 19972
rect 14875 19941 14887 19944
rect 14829 19935 14887 19941
rect 16025 19941 16037 19944
rect 16071 19941 16083 19975
rect 16025 19935 16083 19941
rect 12268 19876 12756 19904
rect 12268 19848 12296 19876
rect 12250 19796 12256 19848
rect 12308 19796 12314 19848
rect 12728 19845 12756 19876
rect 14458 19864 14464 19916
rect 14516 19864 14522 19916
rect 16666 19904 16672 19916
rect 15396 19876 16672 19904
rect 15396 19845 15424 19876
rect 16666 19864 16672 19876
rect 16724 19864 16730 19916
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12713 19839 12771 19845
rect 12575 19808 12609 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12713 19805 12725 19839
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 12544 19768 12572 19799
rect 12802 19768 12808 19780
rect 12176 19740 12808 19768
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 11054 19700 11060 19712
rect 9968 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19700 11118 19712
rect 11149 19703 11207 19709
rect 11149 19700 11161 19703
rect 11112 19672 11161 19700
rect 11112 19660 11118 19672
rect 11149 19669 11161 19672
rect 11195 19669 11207 19703
rect 11149 19663 11207 19669
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 13722 19700 13728 19712
rect 12943 19672 13728 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 14660 19700 14688 19799
rect 15562 19796 15568 19848
rect 15620 19796 15626 19848
rect 15746 19796 15752 19848
rect 15804 19796 15810 19848
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15896 19808 15945 19836
rect 15896 19796 15902 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16206 19796 16212 19848
rect 16264 19796 16270 19848
rect 16390 19796 16396 19848
rect 16448 19836 16454 19848
rect 16868 19845 16896 20012
rect 17678 20000 17684 20012
rect 17736 20040 17742 20052
rect 17736 20012 18368 20040
rect 17736 20000 17742 20012
rect 17865 19975 17923 19981
rect 17865 19941 17877 19975
rect 17911 19941 17923 19975
rect 17865 19935 17923 19941
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19904 17371 19907
rect 17494 19904 17500 19916
rect 17359 19876 17500 19904
rect 17359 19873 17371 19876
rect 17313 19867 17371 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17880 19904 17908 19935
rect 18340 19904 18368 20012
rect 18414 20000 18420 20052
rect 18472 20000 18478 20052
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 18656 20012 18705 20040
rect 18656 20000 18662 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 19518 19904 19524 19916
rect 17880 19876 18276 19904
rect 18340 19876 19524 19904
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 16448 19808 16865 19836
rect 16448 19796 16454 19808
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 16853 19799 16911 19805
rect 17034 19796 17040 19848
rect 17092 19796 17098 19848
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 17586 19836 17592 19848
rect 17451 19808 17592 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 14918 19728 14924 19780
rect 14976 19728 14982 19780
rect 15473 19771 15531 19777
rect 15473 19737 15485 19771
rect 15519 19768 15531 19771
rect 17420 19768 17448 19799
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 18138 19796 18144 19848
rect 18196 19796 18202 19848
rect 18248 19845 18276 19876
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18782 19796 18788 19848
rect 18840 19796 18846 19848
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 18966 19836 18972 19848
rect 18923 19808 18972 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19208 19808 19257 19836
rect 19208 19796 19214 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 15519 19740 17448 19768
rect 17497 19771 17555 19777
rect 15519 19737 15531 19740
rect 15473 19731 15531 19737
rect 17497 19737 17509 19771
rect 17543 19768 17555 19771
rect 18322 19768 18328 19780
rect 17543 19740 18328 19768
rect 17543 19737 17555 19740
rect 17497 19731 17555 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19521 19771 19579 19777
rect 19521 19737 19533 19771
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 16022 19700 16028 19712
rect 14660 19672 16028 19700
rect 16022 19660 16028 19672
rect 16080 19700 16086 19712
rect 16945 19703 17003 19709
rect 16945 19700 16957 19703
rect 16080 19672 16957 19700
rect 16080 19660 16086 19672
rect 16945 19669 16957 19672
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18046 19700 18052 19712
rect 18003 19672 18052 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 19061 19703 19119 19709
rect 19061 19669 19073 19703
rect 19107 19700 19119 19703
rect 19536 19700 19564 19731
rect 19978 19728 19984 19780
rect 20036 19728 20042 19780
rect 19107 19672 19564 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 20990 19660 20996 19712
rect 21048 19660 21054 19712
rect 1104 19610 26864 19632
rect 1104 19558 4829 19610
rect 4881 19558 4893 19610
rect 4945 19558 4957 19610
rect 5009 19558 5021 19610
rect 5073 19558 5085 19610
rect 5137 19558 11268 19610
rect 11320 19558 11332 19610
rect 11384 19558 11396 19610
rect 11448 19558 11460 19610
rect 11512 19558 11524 19610
rect 11576 19558 17707 19610
rect 17759 19558 17771 19610
rect 17823 19558 17835 19610
rect 17887 19558 17899 19610
rect 17951 19558 17963 19610
rect 18015 19558 24146 19610
rect 24198 19558 24210 19610
rect 24262 19558 24274 19610
rect 24326 19558 24338 19610
rect 24390 19558 24402 19610
rect 24454 19558 26864 19610
rect 1104 19536 26864 19558
rect 2866 19496 2872 19508
rect 2746 19468 2872 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2746 19428 2774 19468
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 3335 19499 3393 19505
rect 3335 19496 3347 19499
rect 2976 19468 3347 19496
rect 2976 19428 3004 19468
rect 3335 19465 3347 19468
rect 3381 19465 3393 19499
rect 3335 19459 3393 19465
rect 3421 19499 3479 19505
rect 3421 19465 3433 19499
rect 3467 19496 3479 19499
rect 3467 19468 3648 19496
rect 3467 19465 3479 19468
rect 3421 19459 3479 19465
rect 3620 19428 3648 19468
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 5350 19496 5356 19508
rect 4212 19468 5356 19496
rect 4212 19456 4218 19468
rect 5350 19456 5356 19468
rect 5408 19496 5414 19508
rect 5408 19468 5948 19496
rect 5408 19456 5414 19468
rect 3878 19428 3884 19440
rect 2547 19400 2774 19428
rect 2884 19400 3004 19428
rect 3068 19400 3556 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2406 19320 2412 19372
rect 2464 19320 2470 19372
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2884 19360 2912 19400
rect 3068 19369 3096 19400
rect 3528 19372 3556 19400
rect 3620 19400 3884 19428
rect 2823 19332 2912 19360
rect 2961 19363 3019 19369
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2961 19329 2973 19363
rect 3007 19329 3019 19363
rect 2961 19323 3019 19329
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 3053 19323 3111 19329
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19360 3295 19363
rect 3326 19360 3332 19372
rect 3283 19332 3332 19360
rect 3283 19329 3295 19332
rect 3237 19323 3295 19329
rect 2976 19224 3004 19323
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 3510 19320 3516 19372
rect 3568 19320 3574 19372
rect 3620 19369 3648 19400
rect 3878 19388 3884 19400
rect 3936 19428 3942 19440
rect 5261 19431 5319 19437
rect 3936 19400 5212 19428
rect 3936 19388 3942 19400
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4154 19360 4160 19372
rect 3835 19332 4160 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 4617 19363 4675 19369
rect 4617 19360 4629 19363
rect 4580 19332 4629 19360
rect 4580 19320 4586 19332
rect 4617 19329 4629 19332
rect 4663 19329 4675 19363
rect 5077 19363 5135 19369
rect 5077 19360 5089 19363
rect 4617 19323 4675 19329
rect 4908 19332 5089 19360
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3697 19295 3755 19301
rect 3697 19292 3709 19295
rect 3200 19264 3709 19292
rect 3200 19252 3206 19264
rect 3697 19261 3709 19264
rect 3743 19261 3755 19295
rect 3697 19255 3755 19261
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19292 4767 19295
rect 4798 19292 4804 19304
rect 4755 19264 4804 19292
rect 4755 19261 4767 19264
rect 4709 19255 4767 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 3160 19224 3188 19252
rect 2976 19196 3188 19224
rect 3326 19184 3332 19236
rect 3384 19224 3390 19236
rect 4062 19224 4068 19236
rect 3384 19196 4068 19224
rect 3384 19184 3390 19196
rect 4062 19184 4068 19196
rect 4120 19224 4126 19236
rect 4908 19224 4936 19332
rect 5077 19329 5089 19332
rect 5123 19329 5135 19363
rect 5184 19360 5212 19400
rect 5261 19397 5273 19431
rect 5307 19428 5319 19431
rect 5307 19400 5580 19428
rect 5307 19397 5319 19400
rect 5261 19391 5319 19397
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 5184 19332 5365 19360
rect 5077 19323 5135 19329
rect 5353 19329 5365 19332
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 5445 19363 5503 19369
rect 5445 19329 5457 19363
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19292 5043 19295
rect 5460 19292 5488 19323
rect 5031 19264 5488 19292
rect 5031 19261 5043 19264
rect 4985 19255 5043 19261
rect 4120 19196 4936 19224
rect 4120 19184 4126 19196
rect 2774 19116 2780 19168
rect 2832 19116 2838 19168
rect 5552 19156 5580 19400
rect 5718 19320 5724 19372
rect 5776 19320 5782 19372
rect 5920 19369 5948 19468
rect 9398 19456 9404 19508
rect 9456 19496 9462 19508
rect 10321 19499 10379 19505
rect 10321 19496 10333 19499
rect 9456 19468 10333 19496
rect 9456 19456 9462 19468
rect 10321 19465 10333 19468
rect 10367 19465 10379 19499
rect 10321 19459 10379 19465
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 10594 19496 10600 19508
rect 10468 19468 10600 19496
rect 10468 19456 10474 19468
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 11149 19499 11207 19505
rect 11149 19465 11161 19499
rect 11195 19465 11207 19499
rect 11149 19459 11207 19465
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 11164 19428 11192 19459
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11664 19468 11713 19496
rect 11664 19456 11670 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 16482 19496 16488 19508
rect 14783 19468 16488 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 16482 19456 16488 19468
rect 16540 19496 16546 19508
rect 16540 19468 16712 19496
rect 16540 19456 16546 19468
rect 6972 19400 7130 19428
rect 9416 19400 11192 19428
rect 6972 19388 6978 19400
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 6270 19320 6276 19372
rect 6328 19360 6334 19372
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6328 19332 6377 19360
rect 6328 19320 6334 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 8754 19320 8760 19372
rect 8812 19320 8818 19372
rect 9214 19320 9220 19372
rect 9272 19360 9278 19372
rect 9416 19369 9444 19400
rect 13722 19388 13728 19440
rect 13780 19388 13786 19440
rect 15749 19431 15807 19437
rect 15749 19397 15761 19431
rect 15795 19428 15807 19431
rect 16574 19428 16580 19440
rect 15795 19400 16580 19428
rect 15795 19397 15807 19400
rect 15749 19391 15807 19397
rect 16574 19388 16580 19400
rect 16632 19388 16638 19440
rect 16684 19437 16712 19468
rect 16942 19456 16948 19508
rect 17000 19496 17006 19508
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 17000 19468 17049 19496
rect 17000 19456 17006 19468
rect 17037 19465 17049 19468
rect 17083 19465 17095 19499
rect 19150 19496 19156 19508
rect 17037 19459 17095 19465
rect 17328 19468 19156 19496
rect 16669 19431 16727 19437
rect 16669 19397 16681 19431
rect 16715 19397 16727 19431
rect 16669 19391 16727 19397
rect 16758 19388 16764 19440
rect 16816 19428 16822 19440
rect 17328 19428 17356 19468
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 20901 19499 20959 19505
rect 20901 19496 20913 19499
rect 19576 19468 20913 19496
rect 19576 19456 19582 19468
rect 20901 19465 20913 19468
rect 20947 19465 20959 19499
rect 20901 19459 20959 19465
rect 18874 19428 18880 19440
rect 16816 19400 17356 19428
rect 18814 19400 18880 19428
rect 16816 19388 16822 19400
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9272 19332 9413 19360
rect 9272 19320 9278 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9953 19363 10011 19369
rect 9953 19360 9965 19363
rect 9640 19332 9965 19360
rect 9640 19320 9646 19332
rect 9953 19329 9965 19332
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 10042 19320 10048 19372
rect 10100 19360 10106 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10100 19332 10517 19360
rect 10100 19320 10106 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10652 19332 10977 19360
rect 10652 19320 10658 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 11054 19320 11060 19372
rect 11112 19320 11118 19372
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 11241 19363 11299 19369
rect 11241 19360 11253 19363
rect 11204 19332 11253 19360
rect 11204 19320 11210 19332
rect 11241 19329 11253 19332
rect 11287 19329 11299 19363
rect 11241 19323 11299 19329
rect 11790 19320 11796 19372
rect 11848 19360 11854 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 11848 19332 12173 19360
rect 11848 19320 11854 19332
rect 12161 19329 12173 19332
rect 12207 19360 12219 19363
rect 12526 19360 12532 19372
rect 12207 19332 12532 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16209 19363 16267 19369
rect 16209 19329 16221 19363
rect 16255 19360 16267 19363
rect 16255 19332 16436 19360
rect 16255 19329 16267 19332
rect 16209 19323 16267 19329
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 5644 19264 6653 19292
rect 5644 19233 5672 19264
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 6730 19252 6736 19304
rect 6788 19292 6794 19304
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 6788 19264 8401 19292
rect 6788 19252 6794 19264
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 10870 19292 10876 19304
rect 10827 19264 10876 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 5629 19227 5687 19233
rect 5629 19193 5641 19227
rect 5675 19193 5687 19227
rect 5629 19187 5687 19193
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10597 19227 10655 19233
rect 10597 19224 10609 19227
rect 10284 19196 10609 19224
rect 10284 19184 10290 19196
rect 10597 19193 10609 19196
rect 10643 19193 10655 19227
rect 10704 19224 10732 19255
rect 10870 19252 10876 19264
rect 10928 19292 10934 19304
rect 11698 19292 11704 19304
rect 10928 19264 11704 19292
rect 10928 19252 10934 19264
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 16132 19292 16160 19323
rect 16408 19292 16436 19332
rect 16482 19320 16488 19372
rect 16540 19320 16546 19372
rect 17328 19369 17356 19400
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 19168 19369 19196 19456
rect 20438 19388 20444 19440
rect 20496 19388 20502 19440
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 16758 19292 16764 19304
rect 16132 19264 16252 19292
rect 16408 19264 16764 19292
rect 11054 19224 11060 19236
rect 10704 19196 11060 19224
rect 10597 19187 10655 19193
rect 11054 19184 11060 19196
rect 11112 19224 11118 19236
rect 11882 19224 11888 19236
rect 11112 19196 11888 19224
rect 11112 19184 11118 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 13909 19227 13967 19233
rect 13909 19193 13921 19227
rect 13955 19224 13967 19227
rect 15470 19224 15476 19236
rect 13955 19196 15476 19224
rect 13955 19193 13967 19196
rect 13909 19187 13967 19193
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 15565 19227 15623 19233
rect 15565 19193 15577 19227
rect 15611 19224 15623 19227
rect 15930 19224 15936 19236
rect 15611 19196 15936 19224
rect 15611 19193 15623 19196
rect 15565 19187 15623 19193
rect 15930 19184 15936 19196
rect 15988 19184 15994 19236
rect 16224 19224 16252 19264
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 16390 19224 16396 19236
rect 16224 19196 16396 19224
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 16868 19168 16896 19323
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 18046 19292 18052 19304
rect 17635 19264 18052 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19292 19487 19295
rect 20070 19292 20076 19304
rect 19475 19264 20076 19292
rect 19475 19261 19487 19264
rect 19429 19255 19487 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 5552 19128 6101 19156
rect 6089 19125 6101 19128
rect 6135 19125 6147 19159
rect 6089 19119 6147 19125
rect 12069 19159 12127 19165
rect 12069 19125 12081 19159
rect 12115 19156 12127 19159
rect 12802 19156 12808 19168
rect 12115 19128 12808 19156
rect 12115 19125 12127 19128
rect 12069 19119 12127 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 16758 19156 16764 19168
rect 14240 19128 16764 19156
rect 14240 19116 14246 19128
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 16850 19116 16856 19168
rect 16908 19156 16914 19168
rect 18598 19156 18604 19168
rect 16908 19128 18604 19156
rect 16908 19116 16914 19128
rect 18598 19116 18604 19128
rect 18656 19156 18662 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 18656 19128 19073 19156
rect 18656 19116 18662 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19061 19119 19119 19125
rect 1104 19066 26864 19088
rect 1104 19014 4169 19066
rect 4221 19014 4233 19066
rect 4285 19014 4297 19066
rect 4349 19014 4361 19066
rect 4413 19014 4425 19066
rect 4477 19014 10608 19066
rect 10660 19014 10672 19066
rect 10724 19014 10736 19066
rect 10788 19014 10800 19066
rect 10852 19014 10864 19066
rect 10916 19014 17047 19066
rect 17099 19014 17111 19066
rect 17163 19014 17175 19066
rect 17227 19014 17239 19066
rect 17291 19014 17303 19066
rect 17355 19014 23486 19066
rect 23538 19014 23550 19066
rect 23602 19014 23614 19066
rect 23666 19014 23678 19066
rect 23730 19014 23742 19066
rect 23794 19014 26864 19066
rect 1104 18992 26864 19014
rect 5077 18955 5135 18961
rect 5077 18921 5089 18955
rect 5123 18952 5135 18955
rect 5718 18952 5724 18964
rect 5123 18924 5724 18952
rect 5123 18921 5135 18924
rect 5077 18915 5135 18921
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6914 18912 6920 18964
rect 6972 18912 6978 18964
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 9585 18955 9643 18961
rect 9585 18952 9597 18955
rect 9088 18924 9597 18952
rect 9088 18912 9094 18924
rect 9585 18921 9597 18924
rect 9631 18921 9643 18955
rect 9585 18915 9643 18921
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 10226 18952 10232 18964
rect 9999 18924 10232 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 10965 18955 11023 18961
rect 10965 18952 10977 18955
rect 10560 18924 10977 18952
rect 10560 18912 10566 18924
rect 10965 18921 10977 18924
rect 11011 18921 11023 18955
rect 10965 18915 11023 18921
rect 12526 18912 12532 18964
rect 12584 18912 12590 18964
rect 15378 18912 15384 18964
rect 15436 18952 15442 18964
rect 15565 18955 15623 18961
rect 15565 18952 15577 18955
rect 15436 18924 15577 18952
rect 15436 18912 15442 18924
rect 15565 18921 15577 18924
rect 15611 18921 15623 18955
rect 15565 18915 15623 18921
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 17310 18952 17316 18964
rect 16264 18924 17316 18952
rect 16264 18912 16270 18924
rect 17310 18912 17316 18924
rect 17368 18952 17374 18964
rect 17957 18955 18015 18961
rect 17368 18924 17540 18952
rect 17368 18912 17374 18924
rect 7098 18884 7104 18896
rect 3988 18856 7104 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 3142 18816 3148 18828
rect 1811 18788 3148 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 3513 18819 3571 18825
rect 3513 18816 3525 18819
rect 3384 18788 3525 18816
rect 3384 18776 3390 18788
rect 3513 18785 3525 18788
rect 3559 18785 3571 18819
rect 3513 18779 3571 18785
rect 1486 18708 1492 18760
rect 1544 18708 1550 18760
rect 2866 18708 2872 18760
rect 2924 18708 2930 18760
rect 3988 18757 4016 18856
rect 4614 18776 4620 18828
rect 4672 18776 4678 18828
rect 4798 18776 4804 18828
rect 4856 18816 4862 18828
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 4856 18788 5273 18816
rect 4856 18776 4862 18788
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4522 18708 4528 18760
rect 4580 18748 4586 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4580 18720 4721 18748
rect 4580 18708 4586 18720
rect 4709 18717 4721 18720
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5166 18708 5172 18760
rect 5224 18708 5230 18760
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5442 18748 5448 18760
rect 5399 18720 5448 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 6840 18757 6868 18856
rect 7098 18844 7104 18856
rect 7156 18844 7162 18896
rect 10410 18844 10416 18896
rect 10468 18884 10474 18896
rect 10689 18887 10747 18893
rect 10689 18884 10701 18887
rect 10468 18856 10701 18884
rect 10468 18844 10474 18856
rect 10689 18853 10701 18856
rect 10735 18853 10747 18887
rect 15930 18884 15936 18896
rect 10689 18847 10747 18853
rect 14384 18856 15936 18884
rect 11054 18816 11060 18828
rect 9784 18788 11060 18816
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8812 18720 9137 18748
rect 8812 18708 8818 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 9214 18708 9220 18760
rect 9272 18708 9278 18760
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18748 9367 18751
rect 9398 18748 9404 18760
rect 9355 18720 9404 18748
rect 9355 18717 9367 18720
rect 9309 18711 9367 18717
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9582 18748 9588 18760
rect 9539 18720 9588 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9784 18757 9812 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 14384 18825 14412 18856
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 16669 18887 16727 18893
rect 16669 18884 16681 18887
rect 16540 18856 16681 18884
rect 16540 18844 16546 18856
rect 16669 18853 16681 18856
rect 16715 18853 16727 18887
rect 16669 18847 16727 18853
rect 16758 18844 16764 18896
rect 16816 18884 16822 18896
rect 16816 18856 17448 18884
rect 16816 18844 16822 18856
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 12943 18788 14105 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 17420 18825 17448 18856
rect 17405 18819 17463 18825
rect 14976 18788 17172 18816
rect 14976 18776 14982 18788
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 10502 18708 10508 18760
rect 10560 18708 10566 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18748 12495 18751
rect 12802 18748 12808 18760
rect 12483 18720 12808 18748
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 5184 18680 5212 18708
rect 5534 18680 5540 18692
rect 5184 18652 5540 18680
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 10796 18680 10824 18711
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 10060 18652 10824 18680
rect 10060 18624 10088 18652
rect 3878 18572 3884 18624
rect 3936 18572 3942 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8352 18584 8953 18612
rect 8352 18572 8358 18584
rect 8941 18581 8953 18584
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 10042 18572 10048 18624
rect 10100 18572 10106 18624
rect 15028 18612 15056 18711
rect 15102 18708 15108 18760
rect 15160 18708 15166 18760
rect 15286 18708 15292 18760
rect 15344 18708 15350 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 15396 18680 15424 18711
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15528 18720 15669 18748
rect 15528 18708 15534 18720
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 15746 18708 15752 18760
rect 15804 18748 15810 18760
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15804 18720 16037 18748
rect 15804 18708 15810 18720
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 15841 18683 15899 18689
rect 15841 18680 15853 18683
rect 15396 18652 15853 18680
rect 15841 18649 15853 18652
rect 15887 18649 15899 18683
rect 15841 18643 15899 18649
rect 15562 18612 15568 18624
rect 15028 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15856 18612 15884 18643
rect 15930 18640 15936 18692
rect 15988 18640 15994 18692
rect 16040 18680 16068 18711
rect 16390 18708 16396 18760
rect 16448 18708 16454 18760
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16850 18748 16856 18760
rect 16623 18720 16856 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 17144 18757 17172 18788
rect 17405 18785 17417 18819
rect 17451 18785 17463 18819
rect 17512 18816 17540 18924
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18138 18952 18144 18964
rect 18003 18924 18144 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 18874 18912 18880 18964
rect 18932 18912 18938 18964
rect 20070 18912 20076 18964
rect 20128 18912 20134 18964
rect 20438 18912 20444 18964
rect 20496 18912 20502 18964
rect 19981 18887 20039 18893
rect 19981 18853 19993 18887
rect 20027 18853 20039 18887
rect 19981 18847 20039 18853
rect 17512 18788 17632 18816
rect 17405 18779 17463 18785
rect 17604 18757 17632 18788
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 18104 18788 18521 18816
rect 18104 18776 18110 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 19429 18819 19487 18825
rect 19429 18785 19441 18819
rect 19475 18816 19487 18819
rect 19794 18816 19800 18828
rect 19475 18788 19800 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 18012 18720 18337 18748
rect 18012 18708 18018 18720
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18598 18748 18604 18760
rect 18463 18720 18604 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 18969 18751 19027 18757
rect 18969 18748 18981 18751
rect 18840 18720 18981 18748
rect 18840 18708 18846 18720
rect 18969 18717 18981 18720
rect 19015 18748 19027 18751
rect 19015 18720 19334 18748
rect 19015 18717 19027 18720
rect 18969 18711 19027 18717
rect 16485 18683 16543 18689
rect 16485 18680 16497 18683
rect 16040 18652 16497 18680
rect 16485 18649 16497 18652
rect 16531 18649 16543 18683
rect 16485 18643 16543 18649
rect 17402 18640 17408 18692
rect 17460 18680 17466 18692
rect 17497 18683 17555 18689
rect 17497 18680 17509 18683
rect 17460 18652 17509 18680
rect 17460 18640 17466 18652
rect 17497 18649 17509 18652
rect 17543 18649 17555 18683
rect 19306 18680 19334 18720
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 19996 18748 20024 18847
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 19996 18720 20269 18748
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 20364 18680 20392 18711
rect 26510 18708 26516 18760
rect 26568 18708 26574 18760
rect 19306 18652 20392 18680
rect 17497 18643 17555 18649
rect 16022 18612 16028 18624
rect 15856 18584 16028 18612
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16206 18572 16212 18624
rect 16264 18572 16270 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17678 18612 17684 18624
rect 17092 18584 17684 18612
rect 17092 18572 17098 18584
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 19426 18612 19432 18624
rect 18380 18584 19432 18612
rect 18380 18572 18386 18584
rect 19426 18572 19432 18584
rect 19484 18612 19490 18624
rect 19613 18615 19671 18621
rect 19613 18612 19625 18615
rect 19484 18584 19625 18612
rect 19484 18572 19490 18584
rect 19613 18581 19625 18584
rect 19659 18612 19671 18615
rect 26329 18615 26387 18621
rect 26329 18612 26341 18615
rect 19659 18584 26341 18612
rect 19659 18581 19671 18584
rect 19613 18575 19671 18581
rect 26329 18581 26341 18584
rect 26375 18581 26387 18615
rect 26329 18575 26387 18581
rect 1104 18522 26864 18544
rect 1104 18470 4829 18522
rect 4881 18470 4893 18522
rect 4945 18470 4957 18522
rect 5009 18470 5021 18522
rect 5073 18470 5085 18522
rect 5137 18470 11268 18522
rect 11320 18470 11332 18522
rect 11384 18470 11396 18522
rect 11448 18470 11460 18522
rect 11512 18470 11524 18522
rect 11576 18470 17707 18522
rect 17759 18470 17771 18522
rect 17823 18470 17835 18522
rect 17887 18470 17899 18522
rect 17951 18470 17963 18522
rect 18015 18470 24146 18522
rect 24198 18470 24210 18522
rect 24262 18470 24274 18522
rect 24326 18470 24338 18522
rect 24390 18470 24402 18522
rect 24454 18470 26864 18522
rect 1104 18448 26864 18470
rect 2774 18408 2780 18420
rect 2746 18368 2780 18408
rect 2832 18368 2838 18420
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18408 4123 18411
rect 5166 18408 5172 18420
rect 4111 18380 5172 18408
rect 4111 18377 4123 18380
rect 4065 18371 4123 18377
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18408 10011 18411
rect 10226 18408 10232 18420
rect 9999 18380 10232 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 14550 18408 14556 18420
rect 13771 18380 14556 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 15102 18368 15108 18420
rect 15160 18408 15166 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 15160 18380 15393 18408
rect 15160 18368 15166 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15562 18408 15568 18420
rect 15381 18371 15439 18377
rect 15488 18380 15568 18408
rect 2593 18343 2651 18349
rect 2593 18309 2605 18343
rect 2639 18340 2651 18343
rect 2746 18340 2774 18368
rect 3878 18340 3884 18352
rect 2639 18312 2774 18340
rect 3818 18312 3884 18340
rect 2639 18309 2651 18312
rect 2593 18303 2651 18309
rect 3878 18300 3884 18312
rect 3936 18300 3942 18352
rect 1486 18232 1492 18284
rect 1544 18272 1550 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 1544 18244 2329 18272
rect 1544 18232 1550 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10226 18272 10232 18284
rect 10091 18244 10232 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 10376 18244 13185 18272
rect 10376 18232 10382 18244
rect 13173 18241 13185 18244
rect 13219 18272 13231 18275
rect 13722 18272 13728 18284
rect 13219 18244 13728 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 13924 18244 14749 18272
rect 10244 18204 10272 18232
rect 12526 18204 12532 18216
rect 10244 18176 12532 18204
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18173 13507 18207
rect 13449 18167 13507 18173
rect 12710 18096 12716 18148
rect 12768 18136 12774 18148
rect 13464 18136 13492 18167
rect 13538 18164 13544 18216
rect 13596 18204 13602 18216
rect 13924 18204 13952 18244
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 13596 18176 13952 18204
rect 13596 18164 13602 18176
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14240 18176 14381 18204
rect 14240 18164 14246 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 14645 18207 14703 18213
rect 14645 18173 14657 18207
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 14660 18136 14688 18167
rect 14826 18164 14832 18216
rect 14884 18164 14890 18216
rect 15488 18204 15516 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 15933 18411 15991 18417
rect 15933 18377 15945 18411
rect 15979 18377 15991 18411
rect 15933 18371 15991 18377
rect 15948 18340 15976 18371
rect 16206 18368 16212 18420
rect 16264 18408 16270 18420
rect 16827 18411 16885 18417
rect 16827 18408 16839 18411
rect 16264 18380 16839 18408
rect 16264 18368 16270 18380
rect 16827 18377 16839 18380
rect 16873 18377 16885 18411
rect 16827 18371 16885 18377
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 17221 18411 17279 18417
rect 17221 18408 17233 18411
rect 17000 18380 17233 18408
rect 17000 18368 17006 18380
rect 17221 18377 17233 18380
rect 17267 18377 17279 18411
rect 17221 18371 17279 18377
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 17368 18380 17632 18408
rect 17368 18368 17374 18380
rect 16096 18343 16154 18349
rect 16096 18340 16108 18343
rect 15580 18312 15976 18340
rect 16040 18312 16108 18340
rect 15580 18281 15608 18312
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16040 18272 16068 18312
rect 16096 18309 16108 18312
rect 16142 18309 16154 18343
rect 16096 18303 16154 18309
rect 16301 18343 16359 18349
rect 16301 18309 16313 18343
rect 16347 18340 16359 18343
rect 17037 18343 17095 18349
rect 16347 18312 16896 18340
rect 16347 18309 16359 18312
rect 16301 18303 16359 18309
rect 16868 18284 16896 18312
rect 17037 18309 17049 18343
rect 17083 18340 17095 18343
rect 17083 18312 17448 18340
rect 17083 18309 17095 18312
rect 17037 18303 17095 18309
rect 15988 18244 16068 18272
rect 15988 18232 15994 18244
rect 16850 18232 16856 18284
rect 16908 18272 16914 18284
rect 17313 18275 17371 18281
rect 17313 18272 17325 18275
rect 16908 18244 17325 18272
rect 16908 18232 16914 18244
rect 17313 18241 17325 18244
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 17420 18204 17448 18312
rect 17604 18281 17632 18380
rect 18966 18368 18972 18420
rect 19024 18368 19030 18420
rect 19337 18411 19395 18417
rect 19337 18377 19349 18411
rect 19383 18408 19395 18411
rect 20990 18408 20996 18420
rect 19383 18380 20996 18408
rect 19383 18377 19395 18380
rect 19337 18371 19395 18377
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18272 17647 18275
rect 19352 18272 19380 18371
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 19426 18300 19432 18352
rect 19484 18300 19490 18352
rect 17635 18244 19380 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 17497 18207 17555 18213
rect 17497 18204 17509 18207
rect 15488 18176 17509 18204
rect 17497 18173 17509 18176
rect 17543 18173 17555 18207
rect 17497 18167 17555 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 15105 18139 15163 18145
rect 15105 18136 15117 18139
rect 12768 18108 13676 18136
rect 14660 18108 15117 18136
rect 12768 18096 12774 18108
rect 13538 18028 13544 18080
rect 13596 18028 13602 18080
rect 13648 18068 13676 18108
rect 15105 18105 15117 18108
rect 15151 18105 15163 18139
rect 15105 18099 15163 18105
rect 16574 18096 16580 18148
rect 16632 18136 16638 18148
rect 16669 18139 16727 18145
rect 16669 18136 16681 18139
rect 16632 18108 16681 18136
rect 16632 18096 16638 18108
rect 16669 18105 16681 18108
rect 16715 18105 16727 18139
rect 16669 18099 16727 18105
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 19536 18136 19564 18167
rect 19392 18108 19564 18136
rect 19392 18096 19398 18108
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 13648 18040 14749 18068
rect 14737 18037 14749 18040
rect 14783 18037 14795 18071
rect 14737 18031 14795 18037
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15930 18068 15936 18080
rect 15528 18040 15936 18068
rect 15528 18028 15534 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16390 18068 16396 18080
rect 16163 18040 16396 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 16850 18028 16856 18080
rect 16908 18028 16914 18080
rect 16942 18028 16948 18080
rect 17000 18068 17006 18080
rect 18322 18068 18328 18080
rect 17000 18040 18328 18068
rect 17000 18028 17006 18040
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 1104 17978 26864 18000
rect 1104 17926 4169 17978
rect 4221 17926 4233 17978
rect 4285 17926 4297 17978
rect 4349 17926 4361 17978
rect 4413 17926 4425 17978
rect 4477 17926 10608 17978
rect 10660 17926 10672 17978
rect 10724 17926 10736 17978
rect 10788 17926 10800 17978
rect 10852 17926 10864 17978
rect 10916 17926 17047 17978
rect 17099 17926 17111 17978
rect 17163 17926 17175 17978
rect 17227 17926 17239 17978
rect 17291 17926 17303 17978
rect 17355 17926 23486 17978
rect 23538 17926 23550 17978
rect 23602 17926 23614 17978
rect 23666 17926 23678 17978
rect 23730 17926 23742 17978
rect 23794 17926 26864 17978
rect 1104 17904 26864 17926
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 6638 17864 6644 17876
rect 3476 17836 6644 17864
rect 3476 17824 3482 17836
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10042 17864 10048 17876
rect 9999 17836 10048 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 11054 17864 11060 17876
rect 10367 17836 11060 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12710 17824 12716 17876
rect 12768 17824 12774 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13538 17864 13544 17876
rect 13495 17836 13544 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 15470 17824 15476 17876
rect 15528 17824 15534 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 16945 17867 17003 17873
rect 16945 17864 16957 17867
rect 16724 17836 16957 17864
rect 16724 17824 16730 17836
rect 16945 17833 16957 17836
rect 16991 17833 17003 17867
rect 16945 17827 17003 17833
rect 10686 17756 10692 17808
rect 10744 17756 10750 17808
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 15746 17796 15752 17808
rect 10928 17768 15752 17796
rect 10928 17756 10934 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 15013 17731 15071 17737
rect 7024 17700 14412 17728
rect 7024 17672 7052 17700
rect 14384 17672 14412 17700
rect 15013 17697 15025 17731
rect 15059 17728 15071 17731
rect 16960 17728 16988 17827
rect 15059 17700 15700 17728
rect 16960 17700 19196 17728
rect 15059 17697 15071 17700
rect 15013 17691 15071 17697
rect 15672 17672 15700 17700
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 992 17632 1409 17660
rect 992 17620 998 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 7006 17620 7012 17672
rect 7064 17620 7070 17672
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9456 17632 9689 17660
rect 9456 17620 9462 17632
rect 9677 17629 9689 17632
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9815 17632 10057 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 10045 17629 10057 17632
rect 10091 17660 10103 17663
rect 10318 17660 10324 17672
rect 10091 17632 10324 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 9692 17592 9720 17623
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 12342 17620 12348 17672
rect 12400 17620 12406 17672
rect 12526 17620 12532 17672
rect 12584 17620 12590 17672
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 10686 17592 10692 17604
rect 9692 17564 10692 17592
rect 10686 17552 10692 17564
rect 10744 17552 10750 17604
rect 11057 17595 11115 17601
rect 11057 17561 11069 17595
rect 11103 17561 11115 17595
rect 12360 17592 12388 17620
rect 13280 17592 13308 17623
rect 12360 17564 13308 17592
rect 11057 17555 11115 17561
rect 1578 17484 1584 17536
rect 1636 17484 1642 17536
rect 5721 17527 5779 17533
rect 5721 17493 5733 17527
rect 5767 17524 5779 17527
rect 6270 17524 6276 17536
rect 5767 17496 6276 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 6270 17484 6276 17496
rect 6328 17484 6334 17536
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 10594 17484 10600 17536
rect 10652 17484 10658 17536
rect 11072 17524 11100 17555
rect 11146 17524 11152 17536
rect 11072 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 13464 17524 13492 17623
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 13998 17660 14004 17672
rect 13780 17632 14004 17660
rect 13780 17620 13786 17632
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 14366 17620 14372 17672
rect 14424 17620 14430 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 13909 17595 13967 17601
rect 13909 17561 13921 17595
rect 13955 17592 13967 17595
rect 15304 17592 15332 17623
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18196 17632 18521 17660
rect 18196 17620 18202 17632
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 19168 17660 19196 17700
rect 21818 17660 21824 17672
rect 19168 17632 21824 17660
rect 18509 17623 18567 17629
rect 21818 17620 21824 17632
rect 21876 17660 21882 17672
rect 22833 17663 22891 17669
rect 22833 17660 22845 17663
rect 21876 17632 22845 17660
rect 21876 17620 21882 17632
rect 22833 17629 22845 17632
rect 22879 17629 22891 17663
rect 22833 17623 22891 17629
rect 13955 17564 15332 17592
rect 15396 17564 21496 17592
rect 13955 17561 13967 17564
rect 13909 17555 13967 17561
rect 15396 17524 15424 17564
rect 13464 17496 15424 17524
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 19058 17524 19064 17536
rect 18739 17496 19064 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 21468 17533 21496 17564
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22566 17595 22624 17601
rect 22566 17592 22578 17595
rect 21692 17564 22578 17592
rect 21692 17552 21698 17564
rect 22566 17561 22578 17564
rect 22612 17561 22624 17595
rect 22566 17555 22624 17561
rect 21453 17527 21511 17533
rect 21453 17493 21465 17527
rect 21499 17493 21511 17527
rect 21453 17487 21511 17493
rect 1104 17434 26864 17456
rect 1104 17382 4829 17434
rect 4881 17382 4893 17434
rect 4945 17382 4957 17434
rect 5009 17382 5021 17434
rect 5073 17382 5085 17434
rect 5137 17382 11268 17434
rect 11320 17382 11332 17434
rect 11384 17382 11396 17434
rect 11448 17382 11460 17434
rect 11512 17382 11524 17434
rect 11576 17382 17707 17434
rect 17759 17382 17771 17434
rect 17823 17382 17835 17434
rect 17887 17382 17899 17434
rect 17951 17382 17963 17434
rect 18015 17382 24146 17434
rect 24198 17382 24210 17434
rect 24262 17382 24274 17434
rect 24326 17382 24338 17434
rect 24390 17382 24402 17434
rect 24454 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 6181 17323 6239 17329
rect 1636 17292 6132 17320
rect 1636 17280 1642 17292
rect 4816 17224 5856 17252
rect 4816 17196 4844 17224
rect 3878 17144 3884 17196
rect 3936 17184 3942 17196
rect 3973 17187 4031 17193
rect 3973 17184 3985 17187
rect 3936 17156 3985 17184
rect 3936 17144 3942 17156
rect 3973 17153 3985 17156
rect 4019 17153 4031 17187
rect 3973 17147 4031 17153
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4203 17156 4752 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 3973 16983 4031 16989
rect 3973 16949 3985 16983
rect 4019 16980 4031 16983
rect 4062 16980 4068 16992
rect 4019 16952 4068 16980
rect 4019 16949 4031 16952
rect 3973 16943 4031 16949
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4724 16980 4752 17156
rect 4798 17144 4804 17196
rect 4856 17144 4862 17196
rect 5074 17193 5080 17196
rect 5068 17147 5080 17193
rect 5074 17144 5080 17147
rect 5132 17144 5138 17196
rect 5828 17116 5856 17224
rect 6104 17184 6132 17292
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 6227 17292 9045 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 12897 17323 12955 17329
rect 12897 17320 12909 17323
rect 11204 17292 12909 17320
rect 11204 17280 11210 17292
rect 12897 17289 12909 17292
rect 12943 17320 12955 17323
rect 14826 17320 14832 17332
rect 12943 17292 14832 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 9766 17252 9772 17264
rect 6748 17224 9772 17252
rect 6748 17184 6776 17224
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 13909 17255 13967 17261
rect 13909 17252 13921 17255
rect 13188 17224 13921 17252
rect 6104 17156 6776 17184
rect 6816 17187 6874 17193
rect 6816 17153 6828 17187
rect 6862 17184 6874 17187
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 6862 17156 8033 17184
rect 6862 17153 6874 17156
rect 6816 17147 6874 17153
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8294 17184 8300 17196
rect 8251 17156 8300 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 13188 17193 13216 17224
rect 13909 17221 13921 17224
rect 13955 17252 13967 17255
rect 14090 17252 14096 17264
rect 13955 17224 14096 17252
rect 13955 17221 13967 17224
rect 13909 17215 13967 17221
rect 14090 17212 14096 17224
rect 14148 17212 14154 17264
rect 14200 17261 14228 17292
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15378 17280 15384 17332
rect 15436 17280 15442 17332
rect 18693 17323 18751 17329
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 19334 17320 19340 17332
rect 18739 17292 19340 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17221 14243 17255
rect 15286 17252 15292 17264
rect 14185 17215 14243 17221
rect 14292 17224 15292 17252
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 10652 17156 11529 17184
rect 10652 17144 10658 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 13722 17184 13728 17196
rect 13495 17156 13728 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 6270 17116 6276 17128
rect 5828 17088 6276 17116
rect 6270 17076 6276 17088
rect 6328 17116 6334 17128
rect 6549 17119 6607 17125
rect 6549 17116 6561 17119
rect 6328 17088 6561 17116
rect 6328 17076 6334 17088
rect 6549 17085 6561 17088
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 8478 17076 8484 17128
rect 8536 17076 8542 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17116 8999 17119
rect 9214 17116 9220 17128
rect 8987 17088 9220 17116
rect 8987 17085 8999 17088
rect 8941 17079 8999 17085
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 8570 17048 8576 17060
rect 7975 17020 8576 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 8864 17048 8892 17079
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9723 17088 9812 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9784 17048 9812 17088
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 10870 17116 10876 17128
rect 10560 17088 10876 17116
rect 10560 17076 10566 17088
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11606 17116 11612 17128
rect 11195 17088 11612 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 14292 17116 14320 17224
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18509 17255 18567 17261
rect 18509 17252 18521 17255
rect 18012 17224 18521 17252
rect 18012 17212 18018 17224
rect 18509 17221 18521 17224
rect 18555 17221 18567 17255
rect 19150 17252 19156 17264
rect 18509 17215 18567 17221
rect 18800 17224 19156 17252
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 14660 17156 14841 17184
rect 14660 17125 14688 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 16758 17184 16764 17196
rect 15979 17156 16764 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 18230 17184 18236 17196
rect 16899 17156 18236 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 18230 17144 18236 17156
rect 18288 17184 18294 17196
rect 18800 17193 18828 17224
rect 19150 17212 19156 17224
rect 19208 17212 19214 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 20286 17224 20729 17252
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20717 17215 20775 17221
rect 18785 17187 18843 17193
rect 18288 17156 18736 17184
rect 18288 17144 18294 17156
rect 12406 17088 14320 17116
rect 14645 17119 14703 17125
rect 10134 17048 10140 17060
rect 8864 17020 10140 17048
rect 10134 17008 10140 17020
rect 10192 17048 10198 17060
rect 11238 17048 11244 17060
rect 10192 17020 11244 17048
rect 10192 17008 10198 17020
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 5534 16980 5540 16992
rect 4724 16952 5540 16980
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 8386 16940 8392 16992
rect 8444 16940 8450 16992
rect 10229 16983 10287 16989
rect 10229 16949 10241 16983
rect 10275 16980 10287 16983
rect 11054 16980 11060 16992
rect 10275 16952 11060 16980
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11701 16983 11759 16989
rect 11701 16949 11713 16983
rect 11747 16980 11759 16983
rect 11790 16980 11796 16992
rect 11747 16952 11796 16980
rect 11747 16949 11759 16952
rect 11701 16943 11759 16949
rect 11790 16940 11796 16952
rect 11848 16980 11854 16992
rect 12406 16980 12434 17088
rect 14645 17085 14657 17119
rect 14691 17085 14703 17119
rect 14645 17079 14703 17085
rect 15654 17076 15660 17128
rect 15712 17076 15718 17128
rect 13541 17051 13599 17057
rect 13541 17048 13553 17051
rect 13096 17020 13553 17048
rect 11848 16952 12434 16980
rect 11848 16940 11854 16952
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13096 16989 13124 17020
rect 13541 17017 13553 17020
rect 13587 17017 13599 17051
rect 13541 17011 13599 17017
rect 13630 17008 13636 17060
rect 13688 17048 13694 17060
rect 14461 17051 14519 17057
rect 14461 17048 14473 17051
rect 13688 17020 14473 17048
rect 13688 17008 13694 17020
rect 14461 17017 14473 17020
rect 14507 17017 14519 17051
rect 14461 17011 14519 17017
rect 15013 17051 15071 17057
rect 15013 17017 15025 17051
rect 15059 17048 15071 17051
rect 15838 17048 15844 17060
rect 15059 17020 15844 17048
rect 15059 17017 15071 17020
rect 15013 17011 15071 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 18141 17051 18199 17057
rect 18141 17017 18153 17051
rect 18187 17048 18199 17051
rect 18322 17048 18328 17060
rect 18187 17020 18328 17048
rect 18187 17017 18199 17020
rect 18141 17011 18199 17017
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 18708 17048 18736 17156
rect 18785 17153 18797 17187
rect 18831 17153 18843 17187
rect 18785 17147 18843 17153
rect 20806 17144 20812 17196
rect 20864 17144 20870 17196
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17184 22891 17187
rect 22922 17184 22928 17196
rect 22879 17156 22928 17184
rect 22879 17153 22891 17156
rect 22833 17147 22891 17153
rect 22922 17144 22928 17156
rect 22980 17144 22986 17196
rect 23014 17144 23020 17196
rect 23072 17144 23078 17196
rect 19058 17076 19064 17128
rect 19116 17076 19122 17128
rect 18782 17048 18788 17060
rect 18708 17020 18788 17048
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12860 16952 13093 16980
rect 12860 16940 12866 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13780 16952 13921 16980
rect 13780 16940 13786 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 14093 16983 14151 16989
rect 14093 16980 14105 16983
rect 14056 16952 14105 16980
rect 14056 16940 14062 16952
rect 14093 16949 14105 16952
rect 14139 16949 14151 16983
rect 14093 16943 14151 16949
rect 15746 16940 15752 16992
rect 15804 16940 15810 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 16761 16983 16819 16989
rect 16761 16980 16773 16983
rect 16724 16952 16773 16980
rect 16724 16940 16730 16952
rect 16761 16949 16773 16952
rect 16807 16949 16819 16983
rect 16761 16943 16819 16949
rect 18230 16940 18236 16992
rect 18288 16980 18294 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18288 16952 18521 16980
rect 18288 16940 18294 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 20533 16983 20591 16989
rect 20533 16980 20545 16983
rect 19300 16952 20545 16980
rect 19300 16940 19306 16952
rect 20533 16949 20545 16952
rect 20579 16949 20591 16983
rect 20533 16943 20591 16949
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 22152 16952 22845 16980
rect 22152 16940 22158 16952
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 1104 16890 26864 16912
rect 1104 16838 4169 16890
rect 4221 16838 4233 16890
rect 4285 16838 4297 16890
rect 4349 16838 4361 16890
rect 4413 16838 4425 16890
rect 4477 16838 10608 16890
rect 10660 16838 10672 16890
rect 10724 16838 10736 16890
rect 10788 16838 10800 16890
rect 10852 16838 10864 16890
rect 10916 16838 17047 16890
rect 17099 16838 17111 16890
rect 17163 16838 17175 16890
rect 17227 16838 17239 16890
rect 17291 16838 17303 16890
rect 17355 16838 23486 16890
rect 23538 16838 23550 16890
rect 23602 16838 23614 16890
rect 23666 16838 23678 16890
rect 23730 16838 23742 16890
rect 23794 16838 26864 16890
rect 1104 16816 26864 16838
rect 4798 16776 4804 16788
rect 1688 16748 4804 16776
rect 1688 16652 1716 16748
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 1670 16640 1676 16652
rect 1544 16612 1676 16640
rect 1544 16600 1550 16612
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 3804 16649 3832 16748
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 5132 16748 5273 16776
rect 5132 16736 5138 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 8294 16776 8300 16788
rect 5592 16748 8300 16776
rect 5592 16736 5598 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8536 16748 8769 16776
rect 8536 16736 8542 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 9769 16779 9827 16785
rect 9272 16748 9720 16776
rect 9272 16736 9278 16748
rect 3789 16643 3847 16649
rect 3789 16609 3801 16643
rect 3835 16609 3847 16643
rect 5552 16640 5580 16736
rect 8570 16708 8576 16720
rect 8220 16680 8576 16708
rect 3789 16603 3847 16609
rect 5460 16612 5580 16640
rect 4062 16581 4068 16584
rect 4056 16535 4068 16581
rect 4120 16572 4126 16584
rect 4120 16544 4156 16572
rect 4062 16532 4068 16535
rect 4120 16532 4126 16544
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5460 16581 5488 16612
rect 6270 16600 6276 16652
rect 6328 16600 6334 16652
rect 8220 16649 8248 16680
rect 8570 16668 8576 16680
rect 8628 16708 8634 16720
rect 9398 16708 9404 16720
rect 8628 16680 9404 16708
rect 8628 16668 8634 16680
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 9692 16708 9720 16748
rect 9769 16745 9781 16779
rect 9815 16776 9827 16779
rect 9858 16776 9864 16788
rect 9815 16748 9864 16776
rect 9815 16745 9827 16748
rect 9769 16739 9827 16745
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10965 16779 11023 16785
rect 10459 16748 10916 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 9692 16680 10364 16708
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 8536 16612 9505 16640
rect 8536 16600 8542 16612
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 9824 16612 10180 16640
rect 9824 16600 9830 16612
rect 5261 16575 5319 16581
rect 5261 16572 5273 16575
rect 5132 16544 5273 16572
rect 5132 16532 5138 16544
rect 5261 16541 5273 16544
rect 5307 16541 5319 16575
rect 5261 16535 5319 16541
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16541 5503 16575
rect 5445 16535 5503 16541
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 10152 16581 10180 16612
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 10336 16572 10364 16680
rect 10888 16640 10916 16748
rect 10965 16745 10977 16779
rect 11011 16776 11023 16779
rect 11238 16776 11244 16788
rect 11011 16748 11244 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 11606 16736 11612 16788
rect 11664 16736 11670 16788
rect 13449 16779 13507 16785
rect 13449 16745 13461 16779
rect 13495 16776 13507 16779
rect 13538 16776 13544 16788
rect 13495 16748 13544 16776
rect 13495 16745 13507 16748
rect 13449 16739 13507 16745
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 17034 16776 17040 16788
rect 15804 16748 17040 16776
rect 15804 16736 15810 16748
rect 17034 16736 17040 16748
rect 17092 16776 17098 16788
rect 17954 16776 17960 16788
rect 17092 16748 17960 16776
rect 17092 16736 17098 16748
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 18509 16779 18567 16785
rect 18509 16776 18521 16779
rect 18472 16748 18521 16776
rect 18472 16736 18478 16748
rect 18509 16745 18521 16748
rect 18555 16776 18567 16779
rect 18690 16776 18696 16788
rect 18555 16748 18696 16776
rect 18555 16745 18567 16748
rect 18509 16739 18567 16745
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 19426 16736 19432 16788
rect 19484 16736 19490 16788
rect 22922 16776 22928 16788
rect 21744 16748 22928 16776
rect 11256 16708 11284 16736
rect 15194 16708 15200 16720
rect 11256 16680 11744 16708
rect 11606 16640 11612 16652
rect 10888 16612 11612 16640
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 10689 16575 10747 16581
rect 10689 16572 10701 16575
rect 10336 16544 10701 16572
rect 10137 16535 10195 16541
rect 10689 16541 10701 16544
rect 10735 16541 10747 16575
rect 11716 16572 11744 16680
rect 12452 16680 15200 16708
rect 12452 16649 12480 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 16853 16711 16911 16717
rect 16853 16708 16865 16711
rect 15856 16680 16865 16708
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 12342 16572 12348 16584
rect 10689 16535 10747 16541
rect 10796 16544 11560 16572
rect 11716 16544 12348 16572
rect 1940 16507 1998 16513
rect 1940 16473 1952 16507
rect 1986 16504 1998 16507
rect 2222 16504 2228 16516
rect 1986 16476 2228 16504
rect 1986 16473 1998 16476
rect 1940 16467 1998 16473
rect 2222 16464 2228 16476
rect 2280 16464 2286 16516
rect 3329 16507 3387 16513
rect 3329 16504 3341 16507
rect 3068 16476 3341 16504
rect 2866 16396 2872 16448
rect 2924 16436 2930 16448
rect 3068 16445 3096 16476
rect 3329 16473 3341 16476
rect 3375 16473 3387 16507
rect 3329 16467 3387 16473
rect 3513 16507 3571 16513
rect 3513 16473 3525 16507
rect 3559 16504 3571 16507
rect 3786 16504 3792 16516
rect 3559 16476 3792 16504
rect 3559 16473 3571 16476
rect 3513 16467 3571 16473
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 6546 16513 6552 16516
rect 6540 16504 6552 16513
rect 6507 16476 6552 16504
rect 6540 16467 6552 16476
rect 6546 16464 6552 16467
rect 6604 16464 6610 16516
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 10796 16504 10824 16544
rect 6696 16476 10824 16504
rect 6696 16464 6702 16476
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 11112 16476 11253 16504
rect 11112 16464 11118 16476
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 11330 16464 11336 16516
rect 11388 16504 11394 16516
rect 11425 16507 11483 16513
rect 11425 16504 11437 16507
rect 11388 16476 11437 16504
rect 11388 16464 11394 16476
rect 11425 16473 11437 16476
rect 11471 16473 11483 16507
rect 11532 16504 11560 16544
rect 12342 16532 12348 16544
rect 12400 16572 12406 16584
rect 12820 16572 12848 16603
rect 14090 16600 14096 16652
rect 14148 16600 14154 16652
rect 12400 16544 12848 16572
rect 12400 16532 12406 16544
rect 12894 16532 12900 16584
rect 12952 16572 12958 16584
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12952 16544 13093 16572
rect 12952 16532 12958 16544
rect 13081 16541 13093 16544
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 15856 16572 15884 16680
rect 16853 16677 16865 16680
rect 16899 16677 16911 16711
rect 17972 16708 18000 16736
rect 18877 16711 18935 16717
rect 18877 16708 18889 16711
rect 17972 16680 18889 16708
rect 16853 16671 16911 16677
rect 18877 16677 18889 16680
rect 18923 16677 18935 16711
rect 18877 16671 18935 16677
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19242 16708 19248 16720
rect 19024 16680 19248 16708
rect 19024 16668 19030 16680
rect 19242 16668 19248 16680
rect 19300 16708 19306 16720
rect 19300 16680 19564 16708
rect 19300 16668 19306 16680
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16632 16612 17141 16640
rect 16632 16600 16638 16612
rect 17129 16609 17141 16612
rect 17175 16640 17187 16643
rect 18414 16640 18420 16652
rect 17175 16612 18420 16640
rect 17175 16609 17187 16612
rect 17129 16603 17187 16609
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18782 16600 18788 16652
rect 18840 16640 18846 16652
rect 19536 16649 19564 16680
rect 19521 16643 19579 16649
rect 18840 16612 19472 16640
rect 18840 16600 18846 16612
rect 14792 16544 15884 16572
rect 14792 16532 14798 16544
rect 16758 16532 16764 16584
rect 16816 16572 16822 16584
rect 17402 16572 17408 16584
rect 16816 16544 17408 16572
rect 16816 16532 16822 16544
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 18230 16572 18236 16584
rect 17543 16544 18236 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 15013 16507 15071 16513
rect 15013 16504 15025 16507
rect 11532 16476 15025 16504
rect 11425 16467 11483 16473
rect 15013 16473 15025 16476
rect 15059 16473 15071 16507
rect 16850 16504 16856 16516
rect 15013 16467 15071 16473
rect 16040 16476 16856 16504
rect 3053 16439 3111 16445
rect 3053 16436 3065 16439
rect 2924 16408 3065 16436
rect 2924 16396 2930 16408
rect 3053 16405 3065 16408
rect 3099 16405 3111 16439
rect 3053 16399 3111 16405
rect 3142 16396 3148 16448
rect 3200 16396 3206 16448
rect 3804 16436 3832 16464
rect 5074 16436 5080 16448
rect 3804 16408 5080 16436
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5166 16396 5172 16448
rect 5224 16396 5230 16448
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7340 16408 7665 16436
rect 7340 16396 7346 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7653 16399 7711 16405
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 7800 16408 8953 16436
rect 7800 16396 7806 16408
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 10962 16436 10968 16448
rect 10643 16408 10968 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11149 16439 11207 16445
rect 11149 16405 11161 16439
rect 11195 16436 11207 16439
rect 11698 16436 11704 16448
rect 11195 16408 11704 16436
rect 11195 16405 11207 16408
rect 11149 16399 11207 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 11882 16396 11888 16448
rect 11940 16396 11946 16448
rect 12250 16396 12256 16448
rect 12308 16396 12314 16448
rect 12342 16396 12348 16448
rect 12400 16436 12406 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12400 16408 13001 16436
rect 12400 16396 12406 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14737 16439 14795 16445
rect 14737 16436 14749 16439
rect 14332 16408 14749 16436
rect 14332 16396 14338 16408
rect 14737 16405 14749 16408
rect 14783 16405 14795 16439
rect 14737 16399 14795 16405
rect 14826 16396 14832 16448
rect 14884 16436 14890 16448
rect 16040 16436 16068 16476
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17512 16504 17540 16535
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18322 16532 18328 16584
rect 18380 16532 18386 16584
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18564 16544 18613 16572
rect 18564 16532 18570 16544
rect 18601 16541 18613 16544
rect 18647 16572 18659 16575
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 18647 16544 18705 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 18693 16541 18705 16544
rect 18739 16572 18751 16575
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18739 16544 19257 16572
rect 18739 16541 18751 16544
rect 18693 16535 18751 16541
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19444 16572 19472 16612
rect 19521 16609 19533 16643
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 19628 16612 20484 16640
rect 19628 16572 19656 16612
rect 20456 16581 20484 16612
rect 21634 16600 21640 16652
rect 21692 16600 21698 16652
rect 19444 16544 19656 16572
rect 20441 16575 20499 16581
rect 19245 16535 19303 16541
rect 20441 16541 20453 16575
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 21358 16532 21364 16584
rect 21416 16572 21422 16584
rect 21744 16581 21772 16748
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 23072 16748 23121 16776
rect 23072 16736 23078 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23109 16739 23167 16745
rect 23842 16708 23848 16720
rect 22756 16680 23848 16708
rect 21545 16575 21603 16581
rect 21545 16572 21557 16575
rect 21416 16544 21557 16572
rect 21416 16532 21422 16544
rect 21545 16541 21557 16544
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 17000 16476 17540 16504
rect 17681 16507 17739 16513
rect 17000 16464 17006 16476
rect 17681 16473 17693 16507
rect 17727 16504 17739 16507
rect 17727 16476 18184 16504
rect 17727 16473 17739 16476
rect 17681 16467 17739 16473
rect 14884 16408 16068 16436
rect 14884 16396 14890 16408
rect 16298 16396 16304 16448
rect 16356 16396 16362 16448
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 17865 16439 17923 16445
rect 17865 16436 17877 16439
rect 17644 16408 17877 16436
rect 17644 16396 17650 16408
rect 17865 16405 17877 16408
rect 17911 16405 17923 16439
rect 17865 16399 17923 16405
rect 18046 16396 18052 16448
rect 18104 16396 18110 16448
rect 18156 16436 18184 16476
rect 21634 16464 21640 16516
rect 21692 16504 21698 16516
rect 21836 16504 21864 16535
rect 22554 16532 22560 16584
rect 22612 16532 22618 16584
rect 22756 16581 22784 16680
rect 23842 16668 23848 16680
rect 23900 16668 23906 16720
rect 23400 16612 23888 16640
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 21692 16476 21864 16504
rect 21692 16464 21698 16476
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 22925 16507 22983 16513
rect 22925 16504 22937 16507
rect 22336 16476 22937 16504
rect 22336 16464 22342 16476
rect 22925 16473 22937 16476
rect 22971 16504 22983 16507
rect 23400 16504 23428 16612
rect 23860 16581 23888 16612
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16574 23903 16575
rect 23891 16546 23925 16574
rect 23891 16541 23903 16546
rect 23845 16535 23903 16541
rect 22971 16476 23428 16504
rect 22971 16473 22983 16476
rect 22925 16467 22983 16473
rect 18322 16436 18328 16448
rect 18156 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 19794 16396 19800 16448
rect 19852 16396 19858 16448
rect 20346 16396 20352 16448
rect 20404 16396 20410 16448
rect 22462 16396 22468 16448
rect 22520 16396 22526 16448
rect 23198 16396 23204 16448
rect 23256 16436 23262 16448
rect 23676 16436 23704 16535
rect 24026 16532 24032 16584
rect 24084 16532 24090 16584
rect 23256 16408 23704 16436
rect 23937 16439 23995 16445
rect 23256 16396 23262 16408
rect 23937 16405 23949 16439
rect 23983 16436 23995 16439
rect 24026 16436 24032 16448
rect 23983 16408 24032 16436
rect 23983 16405 23995 16408
rect 23937 16399 23995 16405
rect 24026 16396 24032 16408
rect 24084 16396 24090 16448
rect 1104 16346 26864 16368
rect 1104 16294 4829 16346
rect 4881 16294 4893 16346
rect 4945 16294 4957 16346
rect 5009 16294 5021 16346
rect 5073 16294 5085 16346
rect 5137 16294 11268 16346
rect 11320 16294 11332 16346
rect 11384 16294 11396 16346
rect 11448 16294 11460 16346
rect 11512 16294 11524 16346
rect 11576 16294 17707 16346
rect 17759 16294 17771 16346
rect 17823 16294 17835 16346
rect 17887 16294 17899 16346
rect 17951 16294 17963 16346
rect 18015 16294 24146 16346
rect 24198 16294 24210 16346
rect 24262 16294 24274 16346
rect 24326 16294 24338 16346
rect 24390 16294 24402 16346
rect 24454 16294 26864 16346
rect 1104 16272 26864 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 1596 16164 1624 16195
rect 6546 16192 6552 16244
rect 6604 16232 6610 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6604 16204 6837 16232
rect 6604 16192 6610 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 8386 16232 8392 16244
rect 6972 16204 8392 16232
rect 6972 16192 6978 16204
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 9858 16192 9864 16244
rect 9916 16192 9922 16244
rect 9950 16192 9956 16244
rect 10008 16192 10014 16244
rect 11882 16232 11888 16244
rect 11072 16204 11888 16232
rect 1918 16167 1976 16173
rect 1918 16164 1930 16167
rect 1596 16136 1930 16164
rect 1918 16133 1930 16136
rect 1964 16133 1976 16167
rect 1918 16127 1976 16133
rect 3881 16167 3939 16173
rect 3881 16133 3893 16167
rect 3927 16164 3939 16167
rect 3970 16164 3976 16176
rect 3927 16136 3976 16164
rect 3927 16133 3939 16136
rect 3881 16127 3939 16133
rect 3970 16124 3976 16136
rect 4028 16164 4034 16176
rect 4028 16136 5856 16164
rect 4028 16124 4034 16136
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 1412 16028 1440 16059
rect 1670 16056 1676 16108
rect 1728 16056 1734 16108
rect 4985 16099 5043 16105
rect 1780 16068 2774 16096
rect 1780 16028 1808 16068
rect 1412 16000 1808 16028
rect 2746 15960 2774 16068
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5166 16096 5172 16108
rect 5031 16068 5172 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 5718 16096 5724 16108
rect 5675 16068 5724 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 5828 16105 5856 16136
rect 6270 16124 6276 16176
rect 6328 16164 6334 16176
rect 7085 16167 7143 16173
rect 6328 16136 6960 16164
rect 6328 16124 6334 16136
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6546 16096 6552 16108
rect 5859 16068 6552 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6932 16096 6960 16136
rect 7085 16133 7097 16167
rect 7131 16164 7143 16167
rect 7190 16164 7196 16176
rect 7131 16136 7196 16164
rect 7131 16133 7143 16136
rect 7085 16127 7143 16133
rect 7190 16124 7196 16136
rect 7248 16124 7254 16176
rect 7282 16124 7288 16176
rect 7340 16124 7346 16176
rect 7374 16124 7380 16176
rect 7432 16164 7438 16176
rect 7432 16136 9674 16164
rect 7432 16124 7438 16136
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 6932 16068 8493 16096
rect 6825 16059 6883 16065
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 6840 16028 6868 16059
rect 8570 16056 8576 16108
rect 8628 16096 8634 16108
rect 8737 16099 8795 16105
rect 8737 16096 8749 16099
rect 8628 16068 8749 16096
rect 8628 16056 8634 16068
rect 8737 16065 8749 16068
rect 8783 16065 8795 16099
rect 9646 16096 9674 16136
rect 11072 16105 11100 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 13817 16235 13875 16241
rect 13817 16201 13829 16235
rect 13863 16232 13875 16235
rect 14090 16232 14096 16244
rect 13863 16204 14096 16232
rect 13863 16201 13875 16204
rect 13817 16195 13875 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 14274 16192 14280 16244
rect 14332 16192 14338 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 14642 16232 14648 16244
rect 14415 16204 14648 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 17954 16232 17960 16244
rect 14752 16204 17960 16232
rect 12342 16164 12348 16176
rect 12084 16136 12348 16164
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 9646 16068 10425 16096
rect 8737 16059 8795 16065
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 7742 16028 7748 16040
rect 6840 16000 7748 16028
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 10428 16028 10456 16059
rect 11330 16056 11336 16108
rect 11388 16056 11394 16108
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16096 11575 16099
rect 11606 16096 11612 16108
rect 11563 16068 11612 16096
rect 11563 16065 11575 16068
rect 11517 16059 11575 16065
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12084 16096 12112 16136
rect 12342 16124 12348 16136
rect 12400 16124 12406 16176
rect 13078 16124 13084 16176
rect 13136 16124 13142 16176
rect 14752 16105 14780 16204
rect 17954 16192 17960 16204
rect 18012 16232 18018 16244
rect 18012 16204 19104 16232
rect 18012 16192 18018 16204
rect 16666 16164 16672 16176
rect 16238 16136 16672 16164
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 16837 16167 16895 16173
rect 16837 16133 16849 16167
rect 16883 16164 16895 16167
rect 16942 16164 16948 16176
rect 16883 16136 16948 16164
rect 16883 16133 16895 16136
rect 16837 16127 16895 16133
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 17034 16124 17040 16176
rect 17092 16124 17098 16176
rect 17586 16124 17592 16176
rect 17644 16124 17650 16176
rect 18322 16164 18328 16176
rect 18064 16136 18328 16164
rect 11716 16068 12112 16096
rect 14737 16099 14795 16105
rect 11716 16028 11744 16068
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 17052 16096 17080 16124
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16632 16068 17141 16096
rect 16632 16056 16638 16068
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17604 16096 17632 16124
rect 18064 16108 18092 16136
rect 18322 16124 18328 16136
rect 18380 16164 18386 16176
rect 18693 16167 18751 16173
rect 18693 16164 18705 16167
rect 18380 16136 18705 16164
rect 18380 16124 18386 16136
rect 18693 16133 18705 16136
rect 18739 16133 18751 16167
rect 18693 16127 18751 16133
rect 19076 16108 19104 16204
rect 23934 16192 23940 16244
rect 23992 16192 23998 16244
rect 20346 16124 20352 16176
rect 20404 16124 20410 16176
rect 21358 16124 21364 16176
rect 21416 16164 21422 16176
rect 22088 16167 22146 16173
rect 21416 16136 21956 16164
rect 21416 16124 21422 16136
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 17604 16068 17785 16096
rect 17313 16059 17371 16065
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 10428 16000 11744 16028
rect 8113 15991 8171 15997
rect 3697 15963 3755 15969
rect 3697 15960 3709 15963
rect 2746 15932 3709 15960
rect 3697 15929 3709 15932
rect 3743 15929 3755 15963
rect 3697 15923 3755 15929
rect 4062 15920 4068 15972
rect 4120 15960 4126 15972
rect 4249 15963 4307 15969
rect 4249 15960 4261 15963
rect 4120 15932 4261 15960
rect 4120 15920 4126 15932
rect 4249 15929 4261 15932
rect 4295 15929 4307 15963
rect 4249 15923 4307 15929
rect 6733 15963 6791 15969
rect 6733 15929 6745 15963
rect 6779 15960 6791 15963
rect 6914 15960 6920 15972
rect 6779 15932 6920 15960
rect 6779 15929 6791 15932
rect 6733 15923 6791 15929
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7282 15920 7288 15972
rect 7340 15960 7346 15972
rect 8128 15960 8156 15991
rect 12066 15988 12072 16040
rect 12124 15988 12130 16040
rect 12342 15988 12348 16040
rect 12400 15988 12406 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14599 16000 14872 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 11701 15963 11759 15969
rect 11701 15960 11713 15963
rect 7340 15932 8156 15960
rect 10152 15932 11713 15960
rect 7340 15920 7346 15932
rect 7760 15904 7788 15932
rect 10152 15904 10180 15932
rect 11701 15929 11713 15932
rect 11747 15929 11759 15963
rect 11701 15923 11759 15929
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3418 15892 3424 15904
rect 3099 15864 3424 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 3602 15852 3608 15904
rect 3660 15892 3666 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 3660 15864 3893 15892
rect 3660 15852 3666 15864
rect 3881 15861 3893 15864
rect 3927 15861 3939 15895
rect 3881 15855 3939 15861
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15892 4399 15895
rect 4522 15892 4528 15904
rect 4387 15864 4528 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5626 15852 5632 15904
rect 5684 15852 5690 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7374 15892 7380 15904
rect 7147 15864 7380 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7561 15895 7619 15901
rect 7561 15861 7573 15895
rect 7607 15892 7619 15895
rect 7650 15892 7656 15904
rect 7607 15864 7656 15892
rect 7607 15861 7619 15864
rect 7561 15855 7619 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 7742 15852 7748 15904
rect 7800 15852 7806 15904
rect 10134 15852 10140 15904
rect 10192 15852 10198 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10560 15864 10885 15892
rect 10560 15852 10566 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 10873 15855 10931 15861
rect 11238 15852 11244 15904
rect 11296 15852 11302 15904
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 14844 15892 14872 16000
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 16758 15988 16764 16040
rect 16816 16028 16822 16040
rect 17328 16028 17356 16059
rect 18046 16056 18052 16108
rect 18104 16056 18110 16108
rect 18230 16056 18236 16108
rect 18288 16056 18294 16108
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18472 16068 18521 16096
rect 18472 16056 18478 16068
rect 18509 16065 18521 16068
rect 18555 16096 18567 16099
rect 18966 16096 18972 16108
rect 18555 16068 18972 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 19058 16056 19064 16108
rect 19116 16056 19122 16108
rect 21818 16056 21824 16108
rect 21876 16056 21882 16108
rect 21928 16096 21956 16136
rect 22088 16133 22100 16167
rect 22134 16164 22146 16167
rect 22462 16164 22468 16176
rect 22134 16136 22468 16164
rect 22134 16133 22146 16136
rect 22088 16127 22146 16133
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 21928 16068 23428 16096
rect 17589 16031 17647 16037
rect 17589 16028 17601 16031
rect 16816 16000 17601 16028
rect 16816 15988 16822 16000
rect 17589 15997 17601 16000
rect 17635 15997 17647 16031
rect 17589 15991 17647 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 18138 16028 18144 16040
rect 18003 16000 18144 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 16669 15963 16727 15969
rect 16669 15960 16681 15963
rect 16040 15932 16681 15960
rect 16040 15892 16068 15932
rect 16669 15929 16681 15932
rect 16715 15929 16727 15963
rect 17402 15960 17408 15972
rect 16669 15923 16727 15929
rect 16776 15932 17408 15960
rect 14844 15864 16068 15892
rect 16485 15895 16543 15901
rect 16485 15861 16497 15895
rect 16531 15892 16543 15895
rect 16776 15892 16804 15932
rect 17402 15920 17408 15932
rect 17460 15920 17466 15972
rect 16531 15864 16804 15892
rect 16531 15861 16543 15864
rect 16485 15855 16543 15861
rect 16850 15852 16856 15904
rect 16908 15852 16914 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 17000 15864 17233 15892
rect 17000 15852 17006 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17604 15892 17632 15991
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 19334 15988 19340 16040
rect 19392 15988 19398 16040
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 20772 16000 20821 16028
rect 20772 15988 20778 16000
rect 20809 15997 20821 16000
rect 20855 16028 20867 16031
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 20855 16000 21557 16028
rect 20855 15997 20867 16000
rect 20809 15991 20867 15997
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 22888 16000 23305 16028
rect 22888 15988 22894 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23400 16028 23428 16068
rect 24026 16056 24032 16108
rect 24084 16056 24090 16108
rect 24578 16096 24584 16108
rect 24320 16068 24584 16096
rect 24320 16037 24348 16068
rect 24578 16056 24584 16068
rect 24636 16096 24642 16108
rect 24949 16099 25007 16105
rect 24949 16096 24961 16099
rect 24636 16068 24961 16096
rect 24636 16056 24642 16068
rect 24949 16065 24961 16068
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 25096 16068 25145 16096
rect 25096 16056 25102 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 24305 16031 24363 16037
rect 24305 16028 24317 16031
rect 23400 16000 24317 16028
rect 23293 15991 23351 15997
rect 24305 15997 24317 16000
rect 24351 15997 24363 16031
rect 24305 15991 24363 15997
rect 24121 15963 24179 15969
rect 24121 15929 24133 15963
rect 24167 15960 24179 15963
rect 24486 15960 24492 15972
rect 24167 15932 24492 15960
rect 24167 15929 24179 15932
rect 24121 15923 24179 15929
rect 24486 15920 24492 15932
rect 24544 15920 24550 15972
rect 18141 15895 18199 15901
rect 18141 15892 18153 15895
rect 17604 15864 18153 15892
rect 17221 15855 17279 15861
rect 18141 15861 18153 15864
rect 18187 15861 18199 15895
rect 18141 15855 18199 15861
rect 20990 15852 20996 15904
rect 21048 15852 21054 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 23198 15892 23204 15904
rect 22612 15864 23204 15892
rect 22612 15852 22618 15864
rect 23198 15852 23204 15864
rect 23256 15852 23262 15904
rect 23382 15852 23388 15904
rect 23440 15892 23446 15904
rect 24029 15895 24087 15901
rect 24029 15892 24041 15895
rect 23440 15864 24041 15892
rect 23440 15852 23446 15864
rect 24029 15861 24041 15864
rect 24075 15861 24087 15895
rect 24029 15855 24087 15861
rect 25130 15852 25136 15904
rect 25188 15852 25194 15904
rect 1104 15802 26864 15824
rect 1104 15750 4169 15802
rect 4221 15750 4233 15802
rect 4285 15750 4297 15802
rect 4349 15750 4361 15802
rect 4413 15750 4425 15802
rect 4477 15750 10608 15802
rect 10660 15750 10672 15802
rect 10724 15750 10736 15802
rect 10788 15750 10800 15802
rect 10852 15750 10864 15802
rect 10916 15750 17047 15802
rect 17099 15750 17111 15802
rect 17163 15750 17175 15802
rect 17227 15750 17239 15802
rect 17291 15750 17303 15802
rect 17355 15750 23486 15802
rect 23538 15750 23550 15802
rect 23602 15750 23614 15802
rect 23666 15750 23678 15802
rect 23730 15750 23742 15802
rect 23794 15750 26864 15802
rect 1104 15728 26864 15750
rect 1578 15648 1584 15700
rect 1636 15648 1642 15700
rect 2222 15648 2228 15700
rect 2280 15688 2286 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2280 15660 2329 15688
rect 2280 15648 2286 15660
rect 2317 15657 2329 15660
rect 2363 15657 2375 15691
rect 2317 15651 2375 15657
rect 2777 15691 2835 15697
rect 2777 15657 2789 15691
rect 2823 15688 2835 15691
rect 3142 15688 3148 15700
rect 2823 15660 3148 15688
rect 2823 15657 2835 15660
rect 2777 15651 2835 15657
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3602 15648 3608 15700
rect 3660 15648 3666 15700
rect 3878 15648 3884 15700
rect 3936 15648 3942 15700
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 8478 15688 8484 15700
rect 7699 15660 8484 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 8570 15648 8576 15700
rect 8628 15648 8634 15700
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11664 15660 11989 15688
rect 11664 15648 11670 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 11977 15651 12035 15657
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 12400 15660 12633 15688
rect 12400 15648 12406 15660
rect 12621 15657 12633 15660
rect 12667 15657 12679 15691
rect 12621 15651 12679 15657
rect 13078 15648 13084 15700
rect 13136 15648 13142 15700
rect 15010 15648 15016 15700
rect 15068 15648 15074 15700
rect 15194 15648 15200 15700
rect 15252 15648 15258 15700
rect 17494 15648 17500 15700
rect 17552 15648 17558 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 19334 15688 19340 15700
rect 19291 15660 19340 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 21634 15648 21640 15700
rect 21692 15648 21698 15700
rect 21818 15648 21824 15700
rect 21876 15688 21882 15700
rect 21876 15660 23336 15688
rect 21876 15648 21882 15660
rect 2866 15580 2872 15632
rect 2924 15620 2930 15632
rect 4614 15620 4620 15632
rect 2924 15592 4620 15620
rect 2924 15580 2930 15592
rect 4614 15580 4620 15592
rect 4672 15620 4678 15632
rect 4672 15592 4844 15620
rect 4672 15580 4678 15592
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 3326 15552 3332 15564
rect 3191 15524 3332 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4062 15552 4068 15564
rect 3936 15524 4068 15552
rect 3936 15512 3942 15524
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 4249 15555 4307 15561
rect 4249 15552 4261 15555
rect 4120 15524 4261 15552
rect 4120 15512 4126 15524
rect 4249 15521 4261 15524
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4816 15561 4844 15592
rect 16850 15580 16856 15632
rect 16908 15620 16914 15632
rect 18046 15620 18052 15632
rect 16908 15592 18052 15620
rect 16908 15580 16914 15592
rect 18046 15580 18052 15592
rect 18104 15620 18110 15632
rect 18322 15620 18328 15632
rect 18104 15592 18328 15620
rect 18104 15580 18110 15592
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 21545 15623 21603 15629
rect 21545 15589 21557 15623
rect 21591 15620 21603 15623
rect 22278 15620 22284 15632
rect 21591 15592 22284 15620
rect 21591 15589 21603 15592
rect 21545 15583 21603 15589
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 4801 15555 4859 15561
rect 4396 15524 4660 15552
rect 4396 15512 4402 15524
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2547 15456 2636 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2608 15357 2636 15456
rect 3418 15444 3424 15496
rect 3476 15444 3482 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4522 15484 4528 15496
rect 4203 15456 4528 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4632 15493 4660 15524
rect 4801 15521 4813 15555
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 9674 15552 9680 15564
rect 6604 15524 9680 15552
rect 6604 15512 6610 15524
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 6270 15484 6276 15496
rect 5215 15456 6276 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 7193 15487 7251 15493
rect 7193 15453 7205 15487
rect 7239 15453 7251 15487
rect 7193 15447 7251 15453
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15385 3295 15419
rect 3237 15379 3295 15385
rect 5436 15419 5494 15425
rect 5436 15385 5448 15419
rect 5482 15416 5494 15419
rect 5626 15416 5632 15428
rect 5482 15388 5632 15416
rect 5482 15385 5494 15388
rect 5436 15379 5494 15385
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15317 2651 15351
rect 2593 15311 2651 15317
rect 2774 15308 2780 15360
rect 2832 15308 2838 15360
rect 3252 15348 3280 15379
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 7208 15416 7236 15447
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7340 15456 7389 15484
rect 7340 15444 7346 15456
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 7742 15444 7748 15496
rect 7800 15444 7806 15496
rect 8404 15493 8432 15524
rect 9674 15512 9680 15524
rect 9732 15552 9738 15564
rect 10042 15552 10048 15564
rect 9732 15524 10048 15552
rect 9732 15512 9738 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 12066 15552 12072 15564
rect 10275 15524 12072 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13906 15552 13912 15564
rect 12820 15524 13912 15552
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 12820 15493 12848 15524
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 16942 15552 16948 15564
rect 15120 15524 16948 15552
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8536 15456 8585 15484
rect 8536 15444 8542 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 12805 15487 12863 15493
rect 12805 15453 12817 15487
rect 12851 15453 12863 15487
rect 12805 15447 12863 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13170 15484 13176 15496
rect 13035 15456 13176 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15120 15493 15148 15524
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 17954 15552 17960 15564
rect 17451 15524 17960 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18782 15512 18788 15564
rect 18840 15552 18846 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 18840 15524 19441 15552
rect 18840 15512 18846 15524
rect 19429 15521 19441 15524
rect 19475 15552 19487 15555
rect 20990 15552 20996 15564
rect 19475 15524 20996 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 23308 15561 23336 15660
rect 23293 15555 23351 15561
rect 23293 15521 23305 15555
rect 23339 15552 23351 15555
rect 24489 15555 24547 15561
rect 24489 15552 24501 15555
rect 23339 15524 24501 15552
rect 23339 15521 23351 15524
rect 23293 15515 23351 15521
rect 24489 15521 24501 15524
rect 24535 15521 24547 15555
rect 24489 15515 24547 15521
rect 14921 15487 14979 15493
rect 14921 15484 14933 15487
rect 14792 15456 14933 15484
rect 14792 15444 14798 15456
rect 14921 15453 14933 15456
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15453 15163 15487
rect 15105 15447 15163 15453
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15528 15456 15669 15484
rect 15528 15444 15534 15456
rect 15657 15453 15669 15456
rect 15703 15484 15715 15487
rect 16298 15484 16304 15496
rect 15703 15456 16304 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 18472 15456 19533 15484
rect 18472 15444 18478 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19886 15444 19892 15496
rect 19944 15444 19950 15496
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15453 20775 15487
rect 20717 15447 20775 15453
rect 6564 15388 7420 15416
rect 3326 15348 3332 15360
rect 3252 15320 3332 15348
rect 3326 15308 3332 15320
rect 3384 15348 3390 15360
rect 6564 15357 6592 15388
rect 7392 15360 7420 15388
rect 10502 15376 10508 15428
rect 10560 15376 10566 15428
rect 11238 15376 11244 15428
rect 11296 15376 11302 15428
rect 15381 15419 15439 15425
rect 15381 15385 15393 15419
rect 15427 15385 15439 15419
rect 15381 15379 15439 15385
rect 15565 15419 15623 15425
rect 15565 15385 15577 15419
rect 15611 15416 15623 15419
rect 16482 15416 16488 15428
rect 15611 15388 16488 15416
rect 15611 15385 15623 15388
rect 15565 15379 15623 15385
rect 4433 15351 4491 15357
rect 4433 15348 4445 15351
rect 3384 15320 4445 15348
rect 3384 15308 3390 15320
rect 4433 15317 4445 15320
rect 4479 15317 4491 15351
rect 4433 15311 4491 15317
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15317 6607 15351
rect 6549 15311 6607 15317
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 7432 15320 7481 15348
rect 7432 15308 7438 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7800 15320 7849 15348
rect 7800 15308 7806 15320
rect 7837 15317 7849 15320
rect 7883 15317 7895 15351
rect 15396 15348 15424 15379
rect 16482 15376 16488 15388
rect 16540 15376 16546 15428
rect 16666 15376 16672 15428
rect 16724 15416 16730 15428
rect 17681 15419 17739 15425
rect 17681 15416 17693 15419
rect 16724 15388 17693 15416
rect 16724 15376 16730 15388
rect 17681 15385 17693 15388
rect 17727 15385 17739 15419
rect 17681 15379 17739 15385
rect 17865 15419 17923 15425
rect 17865 15385 17877 15419
rect 17911 15416 17923 15419
rect 18046 15416 18052 15428
rect 17911 15388 18052 15416
rect 17911 15385 17923 15388
rect 17865 15379 17923 15385
rect 18046 15376 18052 15388
rect 18104 15376 18110 15428
rect 19058 15376 19064 15428
rect 19116 15416 19122 15428
rect 20073 15419 20131 15425
rect 20073 15416 20085 15419
rect 19116 15388 20085 15416
rect 19116 15376 19122 15388
rect 20073 15385 20085 15388
rect 20119 15385 20131 15419
rect 20073 15379 20131 15385
rect 20732 15416 20760 15447
rect 20806 15444 20812 15496
rect 20864 15444 20870 15496
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 22094 15484 22100 15496
rect 21683 15456 22100 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 23037 15487 23095 15493
rect 23037 15453 23049 15487
rect 23083 15484 23095 15487
rect 23382 15484 23388 15496
rect 23083 15456 23388 15484
rect 23083 15453 23095 15456
rect 23037 15447 23095 15453
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 24026 15444 24032 15496
rect 24084 15444 24090 15496
rect 24756 15487 24814 15493
rect 24756 15453 24768 15487
rect 24802 15484 24814 15487
rect 25130 15484 25136 15496
rect 24802 15456 25136 15484
rect 24802 15453 24814 15456
rect 24756 15447 24814 15453
rect 25130 15444 25136 15456
rect 25188 15444 25194 15496
rect 20990 15416 20996 15428
rect 20732 15388 20996 15416
rect 16684 15348 16712 15376
rect 15396 15320 16712 15348
rect 7837 15311 7895 15317
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 18380 15320 19625 15348
rect 18380 15308 18386 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20732 15348 20760 15388
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 21358 15376 21364 15428
rect 21416 15376 21422 15428
rect 19852 15320 20760 15348
rect 19852 15308 19858 15320
rect 20898 15308 20904 15360
rect 20956 15308 20962 15360
rect 21913 15351 21971 15357
rect 21913 15317 21925 15351
rect 21959 15348 21971 15351
rect 22830 15348 22836 15360
rect 21959 15320 22836 15348
rect 21959 15317 21971 15320
rect 21913 15311 21971 15317
rect 22830 15308 22836 15320
rect 22888 15308 22894 15360
rect 22922 15308 22928 15360
rect 22980 15348 22986 15360
rect 23385 15351 23443 15357
rect 23385 15348 23397 15351
rect 22980 15320 23397 15348
rect 22980 15308 22986 15320
rect 23385 15317 23397 15320
rect 23431 15317 23443 15351
rect 23385 15311 23443 15317
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 1104 15258 26864 15280
rect 1104 15206 4829 15258
rect 4881 15206 4893 15258
rect 4945 15206 4957 15258
rect 5009 15206 5021 15258
rect 5073 15206 5085 15258
rect 5137 15206 11268 15258
rect 11320 15206 11332 15258
rect 11384 15206 11396 15258
rect 11448 15206 11460 15258
rect 11512 15206 11524 15258
rect 11576 15206 17707 15258
rect 17759 15206 17771 15258
rect 17823 15206 17835 15258
rect 17887 15206 17899 15258
rect 17951 15206 17963 15258
rect 18015 15206 24146 15258
rect 24198 15206 24210 15258
rect 24262 15206 24274 15258
rect 24326 15206 24338 15258
rect 24390 15206 24402 15258
rect 24454 15206 26864 15258
rect 1104 15184 26864 15206
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 3142 15144 3148 15156
rect 2832 15116 3148 15144
rect 2832 15104 2838 15116
rect 3142 15104 3148 15116
rect 3200 15144 3206 15156
rect 3970 15144 3976 15156
rect 3200 15116 3976 15144
rect 3200 15104 3206 15116
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 5718 15144 5724 15156
rect 5675 15116 5724 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 16574 15144 16580 15156
rect 16224 15116 16580 15144
rect 3050 15036 3056 15088
rect 3108 15036 3114 15088
rect 3269 15079 3327 15085
rect 3269 15045 3281 15079
rect 3315 15076 3327 15079
rect 3786 15076 3792 15088
rect 3315 15048 3792 15076
rect 3315 15045 3327 15048
rect 3269 15039 3327 15045
rect 3786 15036 3792 15048
rect 3844 15076 3850 15088
rect 4062 15076 4068 15088
rect 3844 15048 4068 15076
rect 3844 15036 3850 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 16224 15085 16252 15116
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 16666 15104 16672 15156
rect 16724 15104 16730 15156
rect 18049 15147 18107 15153
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 18230 15144 18236 15156
rect 18095 15116 18236 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 18230 15104 18236 15116
rect 18288 15144 18294 15156
rect 18288 15116 18736 15144
rect 18288 15104 18294 15116
rect 16209 15079 16267 15085
rect 16209 15045 16221 15079
rect 16255 15045 16267 15079
rect 16209 15039 16267 15045
rect 16393 15079 16451 15085
rect 16393 15045 16405 15079
rect 16439 15076 16451 15079
rect 16758 15076 16764 15088
rect 16439 15048 16764 15076
rect 16439 15045 16451 15048
rect 16393 15039 16451 15045
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 15008 6055 15011
rect 6638 15008 6644 15020
rect 6043 14980 6644 15008
rect 6043 14977 6055 14980
rect 5997 14971 6055 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 13078 14968 13084 15020
rect 13136 14968 13142 15020
rect 16224 15008 16252 15039
rect 16758 15036 16764 15048
rect 16816 15036 16822 15088
rect 16942 15036 16948 15088
rect 17000 15076 17006 15088
rect 17865 15079 17923 15085
rect 17865 15076 17877 15079
rect 17000 15048 17877 15076
rect 17000 15036 17006 15048
rect 17865 15045 17877 15048
rect 17911 15076 17923 15079
rect 17911 15048 18644 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16224 14980 16681 15008
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6914 14940 6920 14952
rect 6135 14912 6920 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6914 14900 6920 14912
rect 6972 14940 6978 14952
rect 7282 14940 7288 14952
rect 6972 14912 7288 14940
rect 6972 14900 6978 14912
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 16684 14940 16712 14971
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 18138 15008 18144 15020
rect 17543 14980 18144 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 18138 14968 18144 14980
rect 18196 15008 18202 15020
rect 18196 14980 18552 15008
rect 18196 14968 18202 14980
rect 18414 14940 18420 14952
rect 16684 14912 18420 14940
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 17586 14832 17592 14884
rect 17644 14872 17650 14884
rect 18141 14875 18199 14881
rect 18141 14872 18153 14875
rect 17644 14844 18153 14872
rect 17644 14832 17650 14844
rect 18141 14841 18153 14844
rect 18187 14841 18199 14875
rect 18141 14835 18199 14841
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 2924 14776 3249 14804
rect 2924 14764 2930 14776
rect 3237 14773 3249 14776
rect 3283 14773 3295 14807
rect 3237 14767 3295 14773
rect 3421 14807 3479 14813
rect 3421 14773 3433 14807
rect 3467 14804 3479 14807
rect 3878 14804 3884 14816
rect 3467 14776 3884 14804
rect 3467 14773 3479 14776
rect 3421 14767 3479 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 14792 14776 16037 14804
rect 14792 14764 14798 14776
rect 16025 14773 16037 14776
rect 16071 14773 16083 14807
rect 16025 14767 16083 14773
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 18046 14804 18052 14816
rect 17911 14776 18052 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18322 14764 18328 14816
rect 18380 14764 18386 14816
rect 18524 14804 18552 14980
rect 18616 14940 18644 15048
rect 18708 15017 18736 15116
rect 19886 15104 19892 15156
rect 19944 15104 19950 15156
rect 20990 15104 20996 15156
rect 21048 15104 21054 15156
rect 23753 15147 23811 15153
rect 23753 15113 23765 15147
rect 23799 15144 23811 15147
rect 24486 15144 24492 15156
rect 23799 15116 24492 15144
rect 23799 15113 23811 15116
rect 23753 15107 23811 15113
rect 24486 15104 24492 15116
rect 24544 15104 24550 15156
rect 25038 15104 25044 15156
rect 25096 15144 25102 15156
rect 25133 15147 25191 15153
rect 25133 15144 25145 15147
rect 25096 15116 25145 15144
rect 25096 15104 25102 15116
rect 25133 15113 25145 15116
rect 25179 15113 25191 15147
rect 25133 15107 25191 15113
rect 19904 15076 19932 15104
rect 20898 15076 20904 15088
rect 18892 15048 19932 15076
rect 20746 15048 20904 15076
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 18892 14940 18920 15048
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 23385 15079 23443 15085
rect 23385 15045 23397 15079
rect 23431 15045 23443 15079
rect 23385 15039 23443 15045
rect 23601 15079 23659 15085
rect 23601 15045 23613 15079
rect 23647 15076 23659 15079
rect 24026 15076 24032 15088
rect 23647 15048 24032 15076
rect 23647 15045 23659 15048
rect 23601 15039 23659 15045
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 23400 15008 23428 15039
rect 24026 15036 24032 15048
rect 24084 15036 24090 15088
rect 24504 15076 24532 15104
rect 24504 15048 26188 15076
rect 26160 15017 26188 15048
rect 22888 14980 23428 15008
rect 24765 15011 24823 15017
rect 22888 14968 22894 14980
rect 24765 14977 24777 15011
rect 24811 15008 24823 15011
rect 25409 15011 25467 15017
rect 25409 15008 25421 15011
rect 24811 14980 25421 15008
rect 24811 14977 24823 14980
rect 24765 14971 24823 14977
rect 25409 14977 25421 14980
rect 25455 14977 25467 15011
rect 25409 14971 25467 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 18616 14912 18920 14940
rect 19058 14900 19064 14952
rect 19116 14900 19122 14952
rect 19242 14900 19248 14952
rect 19300 14900 19306 14952
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 24544 14912 24685 14940
rect 24544 14900 24550 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 25038 14900 25044 14952
rect 25096 14940 25102 14952
rect 25866 14940 25872 14952
rect 25096 14912 25872 14940
rect 25096 14900 25102 14912
rect 25866 14900 25872 14912
rect 25924 14940 25930 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25924 14912 25973 14940
rect 25924 14900 25930 14912
rect 25961 14909 25973 14912
rect 26007 14940 26019 14943
rect 26252 14940 26280 14971
rect 26418 14968 26424 15020
rect 26476 14968 26482 15020
rect 26007 14912 26280 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 18708 14844 19288 14872
rect 18708 14804 18736 14844
rect 18524 14776 18736 14804
rect 18874 14764 18880 14816
rect 18932 14764 18938 14816
rect 18969 14807 19027 14813
rect 18969 14773 18981 14807
rect 19015 14804 19027 14807
rect 19150 14804 19156 14816
rect 19015 14776 19156 14804
rect 19015 14773 19027 14776
rect 18969 14767 19027 14773
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 19260 14804 19288 14844
rect 22462 14832 22468 14884
rect 22520 14872 22526 14884
rect 23198 14872 23204 14884
rect 22520 14844 23204 14872
rect 22520 14832 22526 14844
rect 23198 14832 23204 14844
rect 23256 14872 23262 14884
rect 23256 14844 23612 14872
rect 23256 14832 23262 14844
rect 20714 14804 20720 14816
rect 19260 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 22738 14764 22744 14816
rect 22796 14764 22802 14816
rect 23584 14813 23612 14844
rect 24118 14832 24124 14884
rect 24176 14872 24182 14884
rect 24578 14872 24584 14884
rect 24176 14844 24584 14872
rect 24176 14832 24182 14844
rect 24578 14832 24584 14844
rect 24636 14832 24642 14884
rect 23569 14807 23627 14813
rect 23569 14773 23581 14807
rect 23615 14773 23627 14807
rect 23569 14767 23627 14773
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 26421 14807 26479 14813
rect 26421 14804 26433 14807
rect 24268 14776 26433 14804
rect 24268 14764 24274 14776
rect 26421 14773 26433 14776
rect 26467 14773 26479 14807
rect 26421 14767 26479 14773
rect 1104 14714 26864 14736
rect 1104 14662 4169 14714
rect 4221 14662 4233 14714
rect 4285 14662 4297 14714
rect 4349 14662 4361 14714
rect 4413 14662 4425 14714
rect 4477 14662 10608 14714
rect 10660 14662 10672 14714
rect 10724 14662 10736 14714
rect 10788 14662 10800 14714
rect 10852 14662 10864 14714
rect 10916 14662 17047 14714
rect 17099 14662 17111 14714
rect 17163 14662 17175 14714
rect 17227 14662 17239 14714
rect 17291 14662 17303 14714
rect 17355 14662 23486 14714
rect 23538 14662 23550 14714
rect 23602 14662 23614 14714
rect 23666 14662 23678 14714
rect 23730 14662 23742 14714
rect 23794 14662 26864 14714
rect 1104 14640 26864 14662
rect 9306 14560 9312 14612
rect 9364 14560 9370 14612
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 15289 14603 15347 14609
rect 15289 14600 15301 14603
rect 15160 14572 15301 14600
rect 15160 14560 15166 14572
rect 15289 14569 15301 14572
rect 15335 14600 15347 14603
rect 15930 14600 15936 14612
rect 15335 14572 15936 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16574 14560 16580 14612
rect 16632 14560 16638 14612
rect 17218 14560 17224 14612
rect 17276 14560 17282 14612
rect 17678 14600 17684 14612
rect 17420 14572 17684 14600
rect 3326 14532 3332 14544
rect 2976 14504 3332 14532
rect 2976 14473 3004 14504
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 10226 14532 10232 14544
rect 3752 14504 10232 14532
rect 3752 14492 3758 14504
rect 10226 14492 10232 14504
rect 10284 14492 10290 14544
rect 17236 14532 17264 14560
rect 16408 14504 17264 14532
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 3418 14464 3424 14476
rect 3108 14436 3424 14464
rect 3108 14424 3114 14436
rect 3418 14424 3424 14436
rect 3476 14464 3482 14476
rect 8478 14464 8484 14476
rect 3476 14436 4384 14464
rect 3476 14424 3482 14436
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3160 14328 3188 14359
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4154 14356 4160 14408
rect 4212 14356 4218 14408
rect 4246 14356 4252 14408
rect 4304 14356 4310 14408
rect 4356 14405 4384 14436
rect 8404 14436 8484 14464
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4614 14356 4620 14408
rect 4672 14356 4678 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 7190 14396 7196 14408
rect 7147 14368 7196 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 4433 14331 4491 14337
rect 3160 14300 4016 14328
rect 3988 14272 4016 14300
rect 4433 14297 4445 14331
rect 4479 14328 4491 14331
rect 5258 14328 5264 14340
rect 4479 14300 5264 14328
rect 4479 14297 4491 14300
rect 4433 14291 4491 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 6932 14328 6960 14359
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 7742 14356 7748 14408
rect 7800 14356 7806 14408
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 6932 14300 7604 14328
rect 2774 14220 2780 14272
rect 2832 14220 2838 14272
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3384 14232 3801 14260
rect 3384 14220 3390 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 3970 14220 3976 14272
rect 4028 14220 4034 14272
rect 4706 14220 4712 14272
rect 4764 14220 4770 14272
rect 6638 14220 6644 14272
rect 6696 14260 6702 14272
rect 7009 14263 7067 14269
rect 7009 14260 7021 14263
rect 6696 14232 7021 14260
rect 6696 14220 6702 14232
rect 7009 14229 7021 14232
rect 7055 14229 7067 14263
rect 7009 14223 7067 14229
rect 7466 14220 7472 14272
rect 7524 14220 7530 14272
rect 7576 14260 7604 14300
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7852 14328 7880 14359
rect 7926 14356 7932 14408
rect 7984 14396 7990 14408
rect 8404 14405 8432 14436
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 12989 14467 13047 14473
rect 8536 14436 9536 14464
rect 8536 14424 8542 14436
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 7984 14368 8401 14396
rect 7984 14356 7990 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8846 14396 8852 14408
rect 8619 14368 8852 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9398 14356 9404 14408
rect 9456 14356 9462 14408
rect 9508 14405 9536 14436
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 14550 14464 14556 14476
rect 13035 14436 14556 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 16408 14473 16436 14504
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14433 16451 14467
rect 17420 14464 17448 14572
rect 17678 14560 17684 14572
rect 17736 14560 17742 14612
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 18322 14560 18328 14612
rect 18380 14560 18386 14612
rect 18509 14603 18567 14609
rect 18509 14569 18521 14603
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 17788 14504 18368 14532
rect 17788 14473 17816 14504
rect 17773 14467 17831 14473
rect 17773 14464 17785 14467
rect 16393 14427 16451 14433
rect 16684 14436 17448 14464
rect 17512 14436 17785 14464
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9674 14356 9680 14408
rect 9732 14356 9738 14408
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 13688 14368 14657 14396
rect 13688 14356 13694 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14826 14356 14832 14408
rect 14884 14356 14890 14408
rect 14918 14356 14924 14408
rect 14976 14396 14982 14408
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14976 14368 15117 14396
rect 14976 14356 14982 14368
rect 15105 14365 15117 14368
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16574 14396 16580 14408
rect 15795 14368 16580 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16684 14405 16712 14436
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16908 14368 16957 14396
rect 16908 14356 16914 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17313 14399 17371 14405
rect 17313 14365 17325 14399
rect 17359 14396 17371 14399
rect 17402 14396 17408 14408
rect 17359 14368 17408 14396
rect 17359 14365 17371 14368
rect 17313 14359 17371 14365
rect 17402 14356 17408 14368
rect 17460 14396 17466 14408
rect 17512 14396 17540 14436
rect 17773 14433 17785 14436
rect 17819 14433 17831 14467
rect 18046 14464 18052 14476
rect 17773 14427 17831 14433
rect 17880 14436 18052 14464
rect 17880 14405 17908 14436
rect 18046 14424 18052 14436
rect 18104 14464 18110 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18104 14436 18245 14464
rect 18104 14424 18110 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18340 14464 18368 14504
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 18524 14532 18552 14563
rect 18874 14560 18880 14612
rect 18932 14600 18938 14612
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18932 14572 18981 14600
rect 18932 14560 18938 14572
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19518 14600 19524 14612
rect 19383 14572 19524 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 20165 14603 20223 14609
rect 20165 14569 20177 14603
rect 20211 14600 20223 14603
rect 20622 14600 20628 14612
rect 20211 14572 20628 14600
rect 20211 14569 20223 14572
rect 20165 14563 20223 14569
rect 18472 14504 18552 14532
rect 18785 14535 18843 14541
rect 18472 14492 18478 14504
rect 18785 14501 18797 14535
rect 18831 14501 18843 14535
rect 18785 14495 18843 14501
rect 18506 14464 18512 14476
rect 18340 14436 18512 14464
rect 18233 14427 18291 14433
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 18800 14464 18828 14495
rect 19058 14492 19064 14544
rect 19116 14532 19122 14544
rect 19886 14532 19892 14544
rect 19116 14504 19892 14532
rect 19116 14492 19122 14504
rect 19886 14492 19892 14504
rect 19944 14532 19950 14544
rect 20180 14532 20208 14563
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 24854 14600 24860 14612
rect 24136 14572 24860 14600
rect 24136 14541 24164 14572
rect 24854 14560 24860 14572
rect 24912 14560 24918 14612
rect 19944 14504 20208 14532
rect 24121 14535 24179 14541
rect 19944 14492 19950 14504
rect 24121 14501 24133 14535
rect 24167 14501 24179 14535
rect 24121 14495 24179 14501
rect 18966 14464 18972 14476
rect 18800 14436 18972 14464
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 19794 14464 19800 14476
rect 19659 14436 19800 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14464 20039 14467
rect 20714 14464 20720 14476
rect 20027 14436 20720 14464
rect 20027 14433 20039 14436
rect 19981 14427 20039 14433
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14464 23075 14467
rect 23934 14464 23940 14476
rect 23063 14436 23940 14464
rect 23063 14433 23075 14436
rect 23017 14427 23075 14433
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24136 14436 24716 14464
rect 17460 14368 17540 14396
rect 17877 14399 17935 14405
rect 17460 14356 17466 14368
rect 17877 14365 17889 14399
rect 17923 14365 17935 14399
rect 18417 14399 18475 14405
rect 17877 14359 17935 14365
rect 7708 14300 7880 14328
rect 8021 14331 8079 14337
rect 7708 14288 7714 14300
rect 8021 14297 8033 14331
rect 8067 14328 8079 14331
rect 8754 14328 8760 14340
rect 8067 14300 8760 14328
rect 8067 14297 8079 14300
rect 8021 14291 8079 14297
rect 8754 14288 8760 14300
rect 8812 14288 8818 14340
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 12713 14331 12771 14337
rect 12713 14328 12725 14331
rect 12308 14300 12725 14328
rect 12308 14288 12314 14300
rect 12713 14297 12725 14300
rect 12759 14328 12771 14331
rect 14936 14328 14964 14356
rect 12759 14300 14964 14328
rect 12759 14297 12771 14300
rect 12713 14291 12771 14297
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15933 14331 15991 14337
rect 18322 14334 18328 14386
rect 18380 14334 18386 14386
rect 18417 14365 18429 14399
rect 18463 14390 18475 14399
rect 18463 14365 18644 14390
rect 18417 14362 18644 14365
rect 18417 14359 18475 14362
rect 15933 14328 15945 14331
rect 15712 14300 15945 14328
rect 15712 14288 15718 14300
rect 15933 14297 15945 14300
rect 15979 14297 15991 14331
rect 15933 14291 15991 14297
rect 8202 14260 8208 14272
rect 7576 14232 8208 14260
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8720 14232 8953 14260
rect 8720 14220 8726 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9585 14263 9643 14269
rect 9585 14229 9597 14263
rect 9631 14260 9643 14263
rect 9766 14260 9772 14272
rect 9631 14232 9772 14260
rect 9631 14229 9643 14232
rect 9585 14223 9643 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12345 14263 12403 14269
rect 12345 14260 12357 14263
rect 11756 14232 12357 14260
rect 11756 14220 11762 14232
rect 12345 14229 12357 14232
rect 12391 14229 12403 14263
rect 12345 14223 12403 14229
rect 12802 14220 12808 14272
rect 12860 14220 12866 14272
rect 14090 14220 14096 14272
rect 14148 14220 14154 14272
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 15562 14220 15568 14272
rect 15620 14220 15626 14272
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 16761 14263 16819 14269
rect 16761 14260 16773 14263
rect 16724 14232 16773 14260
rect 16724 14220 16730 14232
rect 16761 14229 16773 14232
rect 16807 14229 16819 14263
rect 16761 14223 16819 14229
rect 17494 14220 17500 14272
rect 17552 14220 17558 14272
rect 18616 14260 18644 14362
rect 19058 14356 19064 14408
rect 19116 14356 19122 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19208 14368 19257 14396
rect 19208 14356 19214 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 19444 14328 19472 14359
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 22554 14356 22560 14408
rect 22612 14356 22618 14408
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 22830 14356 22836 14408
rect 22888 14356 22894 14408
rect 22922 14356 22928 14408
rect 22980 14396 22986 14408
rect 23109 14399 23167 14405
rect 23109 14396 23121 14399
rect 22980 14368 23121 14396
rect 22980 14356 22986 14368
rect 23109 14365 23121 14368
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23293 14399 23351 14405
rect 23293 14396 23305 14399
rect 23256 14368 23305 14396
rect 23256 14356 23262 14368
rect 23293 14365 23305 14368
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 24136 14396 24164 14436
rect 23891 14368 24164 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24210 14356 24216 14408
rect 24268 14356 24274 14408
rect 24578 14356 24584 14408
rect 24636 14356 24642 14408
rect 24688 14396 24716 14436
rect 24688 14368 25084 14396
rect 25056 14340 25084 14368
rect 18748 14300 19472 14328
rect 23477 14331 23535 14337
rect 18748 14288 18754 14300
rect 23477 14297 23489 14331
rect 23523 14328 23535 14331
rect 23937 14331 23995 14337
rect 23523 14300 23888 14328
rect 23523 14297 23535 14300
rect 23477 14291 23535 14297
rect 23860 14272 23888 14300
rect 23937 14297 23949 14331
rect 23983 14328 23995 14331
rect 24118 14328 24124 14340
rect 23983 14300 24124 14328
rect 23983 14297 23995 14300
rect 23937 14291 23995 14297
rect 24118 14288 24124 14300
rect 24176 14288 24182 14340
rect 24826 14331 24884 14337
rect 24826 14328 24838 14331
rect 24228 14300 24838 14328
rect 18782 14260 18788 14272
rect 18616 14232 18788 14260
rect 18782 14220 18788 14232
rect 18840 14260 18846 14272
rect 19426 14260 19432 14272
rect 18840 14232 19432 14260
rect 18840 14220 18846 14232
rect 19426 14220 19432 14232
rect 19484 14260 19490 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 19484 14232 19809 14260
rect 19484 14220 19490 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 22186 14220 22192 14272
rect 22244 14260 22250 14272
rect 22373 14263 22431 14269
rect 22373 14260 22385 14263
rect 22244 14232 22385 14260
rect 22244 14220 22250 14232
rect 22373 14229 22385 14232
rect 22419 14229 22431 14263
rect 22373 14223 22431 14229
rect 23750 14220 23756 14272
rect 23808 14220 23814 14272
rect 23842 14220 23848 14272
rect 23900 14220 23906 14272
rect 24228 14269 24256 14300
rect 24826 14297 24838 14300
rect 24872 14297 24884 14331
rect 24826 14291 24884 14297
rect 25038 14288 25044 14340
rect 25096 14288 25102 14340
rect 24213 14263 24271 14269
rect 24213 14229 24225 14263
rect 24259 14229 24271 14263
rect 24213 14223 24271 14229
rect 25958 14220 25964 14272
rect 26016 14220 26022 14272
rect 1104 14170 26864 14192
rect 1104 14118 4829 14170
rect 4881 14118 4893 14170
rect 4945 14118 4957 14170
rect 5009 14118 5021 14170
rect 5073 14118 5085 14170
rect 5137 14118 11268 14170
rect 11320 14118 11332 14170
rect 11384 14118 11396 14170
rect 11448 14118 11460 14170
rect 11512 14118 11524 14170
rect 11576 14118 17707 14170
rect 17759 14118 17771 14170
rect 17823 14118 17835 14170
rect 17887 14118 17899 14170
rect 17951 14118 17963 14170
rect 18015 14118 24146 14170
rect 24198 14118 24210 14170
rect 24262 14118 24274 14170
rect 24326 14118 24338 14170
rect 24390 14118 24402 14170
rect 24454 14118 26864 14170
rect 1104 14096 26864 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 3694 14056 3700 14068
rect 1627 14028 3700 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4246 14056 4252 14068
rect 4019 14028 4252 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 6546 14056 6552 14068
rect 6380 14028 6552 14056
rect 2501 13991 2559 13997
rect 2501 13957 2513 13991
rect 2547 13988 2559 13991
rect 3142 13988 3148 14000
rect 2547 13960 3148 13988
rect 2547 13957 2559 13960
rect 2501 13951 2559 13957
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 6380 13997 6408 14028
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6733 14059 6791 14065
rect 6733 14025 6745 14059
rect 6779 14056 6791 14059
rect 6914 14056 6920 14068
rect 6779 14028 6920 14056
rect 6779 14025 6791 14028
rect 6733 14019 6791 14025
rect 6365 13991 6423 13997
rect 6365 13957 6377 13991
rect 6411 13957 6423 13991
rect 6748 13988 6776 14019
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7190 14016 7196 14068
rect 7248 14016 7254 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8536 14028 8677 14056
rect 8536 14016 8542 14028
rect 8665 14025 8677 14028
rect 8711 14025 8723 14059
rect 8665 14019 8723 14025
rect 9674 14016 9680 14068
rect 9732 14016 9738 14068
rect 13630 14016 13636 14068
rect 13688 14016 13694 14068
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 14550 14016 14556 14068
rect 14608 14016 14614 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15355 14059 15413 14065
rect 15355 14056 15367 14059
rect 14976 14028 15367 14056
rect 14976 14016 14982 14028
rect 15355 14025 15367 14028
rect 15401 14025 15413 14059
rect 18138 14056 18144 14068
rect 15355 14019 15413 14025
rect 17420 14028 18144 14056
rect 6365 13951 6423 13957
rect 6564 13960 6776 13988
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 4062 13920 4068 13932
rect 2915 13892 4068 13920
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4982 13880 4988 13932
rect 5040 13880 5046 13932
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 6564 13929 6592 13960
rect 6871 13957 6929 13963
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 5224 13892 5365 13920
rect 5224 13880 5230 13892
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6871 13923 6883 13957
rect 6917 13923 6929 13957
rect 7098 13948 7104 14000
rect 7156 13948 7162 14000
rect 7926 13988 7932 14000
rect 7392 13960 7932 13988
rect 6871 13920 6929 13923
rect 7392 13920 7420 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8260 13960 9904 13988
rect 8260 13948 8266 13960
rect 6871 13917 7420 13920
rect 6886 13892 7420 13917
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 8113 13923 8171 13929
rect 8113 13920 8125 13923
rect 7524 13892 8125 13920
rect 7524 13880 7530 13892
rect 8113 13889 8125 13892
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 3476 13824 4169 13852
rect 3476 13812 3482 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 5184 13852 5212 13880
rect 4157 13815 4215 13821
rect 4264 13824 5212 13852
rect 5261 13855 5319 13861
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4264 13784 4292 13824
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5534 13852 5540 13864
rect 5307 13824 5540 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7156 13824 7757 13852
rect 7156 13812 7162 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 8312 13852 8340 13883
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13920 8539 13923
rect 8570 13920 8576 13932
rect 8527 13892 8576 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 9766 13880 9772 13932
rect 9824 13880 9830 13932
rect 9876 13929 9904 13960
rect 10042 13948 10048 14000
rect 10100 13948 10106 14000
rect 12066 13988 12072 14000
rect 11900 13960 12072 13988
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 11606 13920 11612 13932
rect 10827 13892 11612 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 11900 13929 11928 13960
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 13538 13988 13544 14000
rect 13386 13960 13544 13988
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 14185 13991 14243 13997
rect 14185 13957 14197 13991
rect 14231 13988 14243 13991
rect 15010 13988 15016 14000
rect 14231 13960 15016 13988
rect 14231 13957 14243 13960
rect 14185 13951 14243 13957
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 15565 13991 15623 13997
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 17420 13988 17448 14028
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 18690 14056 18696 14068
rect 18279 14028 18696 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 22554 14016 22560 14068
rect 22612 14016 22618 14068
rect 22646 14016 22652 14068
rect 22704 14056 22710 14068
rect 22925 14059 22983 14065
rect 22925 14056 22937 14059
rect 22704 14028 22937 14056
rect 22704 14016 22710 14028
rect 22925 14025 22937 14028
rect 22971 14025 22983 14059
rect 22925 14019 22983 14025
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25314 14056 25320 14068
rect 24912 14028 25320 14056
rect 24912 14016 24918 14028
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 26418 14016 26424 14068
rect 26476 14016 26482 14068
rect 15611 13960 17448 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15105 13923 15163 13929
rect 15105 13920 15117 13923
rect 14976 13892 15117 13920
rect 14976 13880 14982 13892
rect 15105 13889 15117 13892
rect 15151 13920 15163 13923
rect 15580 13920 15608 13951
rect 17328 13929 17356 13960
rect 18322 13948 18328 14000
rect 18380 13948 18386 14000
rect 22572 13988 22600 14016
rect 22833 13991 22891 13997
rect 22833 13988 22845 13991
rect 22572 13960 22845 13988
rect 22833 13957 22845 13960
rect 22879 13957 22891 13991
rect 23201 13991 23259 13997
rect 23201 13988 23213 13991
rect 22833 13951 22891 13957
rect 22940 13960 23213 13988
rect 15151 13892 15608 13920
rect 17313 13923 17371 13929
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 17313 13889 17325 13923
rect 17359 13889 17371 13923
rect 17313 13883 17371 13889
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13920 17647 13923
rect 18340 13920 18368 13948
rect 18598 13920 18604 13932
rect 17635 13892 18604 13920
rect 17635 13889 17647 13892
rect 17589 13883 17647 13889
rect 8312 13824 8432 13852
rect 7745 13815 7803 13821
rect 4028 13756 4292 13784
rect 4028 13744 4034 13756
rect 4522 13744 4528 13796
rect 4580 13744 4586 13796
rect 7558 13744 7564 13796
rect 7616 13784 7622 13796
rect 8404 13784 8432 13824
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8904 13824 9045 13852
rect 8904 13812 8910 13824
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 12158 13812 12164 13864
rect 12216 13812 12222 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15010 13852 15016 13864
rect 14875 13824 15016 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 9122 13784 9128 13796
rect 7616 13756 9128 13784
rect 7616 13744 7622 13756
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 13170 13744 13176 13796
rect 13228 13784 13234 13796
rect 13725 13787 13783 13793
rect 13725 13784 13737 13787
rect 13228 13756 13737 13784
rect 13228 13744 13234 13756
rect 13725 13753 13737 13756
rect 13771 13753 13783 13787
rect 14384 13784 14412 13815
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 17420 13852 17448 13883
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22370 13880 22376 13932
rect 22428 13880 22434 13932
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13920 22615 13923
rect 22738 13920 22744 13932
rect 22603 13892 22744 13920
rect 22603 13889 22615 13892
rect 22557 13883 22615 13889
rect 17494 13852 17500 13864
rect 17420 13824 17500 13852
rect 15197 13787 15255 13793
rect 15197 13784 15209 13787
rect 14384 13756 15209 13784
rect 13725 13747 13783 13753
rect 15197 13753 15209 13756
rect 15243 13753 15255 13787
rect 17420 13784 17448 13824
rect 17494 13812 17500 13824
rect 17552 13852 17558 13864
rect 18322 13852 18328 13864
rect 17552 13824 18328 13852
rect 17552 13812 17558 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 19794 13852 19800 13864
rect 18555 13824 19800 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 15197 13747 15255 13753
rect 15304 13756 17448 13784
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 1728 13688 2329 13716
rect 1728 13676 1734 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2317 13679 2375 13685
rect 2501 13719 2559 13725
rect 2501 13685 2513 13719
rect 2547 13716 2559 13719
rect 2774 13716 2780 13728
rect 2547 13688 2780 13716
rect 2547 13685 2559 13688
rect 2501 13679 2559 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 4614 13676 4620 13728
rect 4672 13676 4678 13728
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 4801 13719 4859 13725
rect 4801 13716 4813 13719
rect 4764 13688 4813 13716
rect 4764 13676 4770 13688
rect 4801 13685 4813 13688
rect 4847 13685 4859 13719
rect 4801 13679 4859 13685
rect 5166 13676 5172 13728
rect 5224 13676 5230 13728
rect 5442 13676 5448 13728
rect 5500 13676 5506 13728
rect 6454 13676 6460 13728
rect 6512 13676 6518 13728
rect 6917 13719 6975 13725
rect 6917 13685 6929 13719
rect 6963 13716 6975 13719
rect 7834 13716 7840 13728
rect 6963 13688 7840 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 7834 13676 7840 13688
rect 7892 13716 7898 13728
rect 8846 13716 8852 13728
rect 7892 13688 8852 13716
rect 7892 13676 7898 13688
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 9953 13719 10011 13725
rect 9953 13685 9965 13719
rect 9999 13716 10011 13719
rect 10042 13716 10048 13728
rect 9999 13688 10048 13716
rect 9999 13685 10011 13688
rect 9953 13679 10011 13685
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 11054 13716 11060 13728
rect 11011 13688 11060 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11517 13719 11575 13725
rect 11517 13716 11529 13719
rect 11204 13688 11529 13716
rect 11204 13676 11210 13688
rect 11517 13685 11529 13688
rect 11563 13685 11575 13719
rect 11517 13679 11575 13685
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 14884 13688 15025 13716
rect 14884 13676 14890 13688
rect 15013 13685 15025 13688
rect 15059 13716 15071 13719
rect 15304 13716 15332 13756
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18524 13784 18552 13815
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22480 13852 22508 13883
rect 22738 13880 22744 13892
rect 22796 13920 22802 13932
rect 22940 13920 22968 13960
rect 23201 13957 23213 13960
rect 23247 13957 23259 13991
rect 23201 13951 23259 13957
rect 24486 13948 24492 14000
rect 24544 13988 24550 14000
rect 25009 13991 25067 13997
rect 25009 13988 25021 13991
rect 24544 13960 25021 13988
rect 24544 13948 24550 13960
rect 25009 13957 25021 13960
rect 25055 13957 25067 13991
rect 25009 13951 25067 13957
rect 25225 13991 25283 13997
rect 25225 13957 25237 13991
rect 25271 13957 25283 13991
rect 25225 13951 25283 13957
rect 22796 13892 22968 13920
rect 22796 13880 22802 13892
rect 23014 13880 23020 13932
rect 23072 13920 23078 13932
rect 23109 13923 23167 13929
rect 23109 13920 23121 13923
rect 23072 13892 23121 13920
rect 23072 13880 23078 13892
rect 23109 13889 23121 13892
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 23290 13880 23296 13932
rect 23348 13880 23354 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23750 13920 23756 13932
rect 23532 13892 23756 13920
rect 23532 13880 23538 13892
rect 23750 13880 23756 13892
rect 23808 13880 23814 13932
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13920 23995 13923
rect 25240 13920 25268 13951
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 23983 13892 25789 13920
rect 23983 13889 23995 13892
rect 23937 13883 23995 13889
rect 25777 13889 25789 13892
rect 25823 13920 25835 13923
rect 25958 13920 25964 13932
rect 25823 13892 25964 13920
rect 25823 13889 25835 13892
rect 25777 13883 25835 13889
rect 25958 13880 25964 13892
rect 26016 13880 26022 13932
rect 22152 13824 22876 13852
rect 22152 13812 22158 13824
rect 18104 13756 18552 13784
rect 22848 13784 22876 13824
rect 22922 13812 22928 13864
rect 22980 13852 22986 13864
rect 23845 13855 23903 13861
rect 23845 13852 23857 13855
rect 22980 13824 23857 13852
rect 22980 13812 22986 13824
rect 23845 13821 23857 13824
rect 23891 13821 23903 13855
rect 23845 13815 23903 13821
rect 24670 13812 24676 13864
rect 24728 13812 24734 13864
rect 23014 13784 23020 13796
rect 22848 13756 23020 13784
rect 18104 13744 18110 13756
rect 23014 13744 23020 13756
rect 23072 13744 23078 13796
rect 15059 13688 15332 13716
rect 15059 13685 15071 13688
rect 15013 13679 15071 13685
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 16942 13716 16948 13728
rect 15436 13688 16948 13716
rect 15436 13676 15442 13688
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 18601 13719 18659 13725
rect 18601 13685 18613 13719
rect 18647 13716 18659 13719
rect 18874 13716 18880 13728
rect 18647 13688 18880 13716
rect 18647 13685 18659 13688
rect 18601 13679 18659 13685
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 24026 13676 24032 13728
rect 24084 13676 24090 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 26864 13648
rect 1104 13574 4169 13626
rect 4221 13574 4233 13626
rect 4285 13574 4297 13626
rect 4349 13574 4361 13626
rect 4413 13574 4425 13626
rect 4477 13574 10608 13626
rect 10660 13574 10672 13626
rect 10724 13574 10736 13626
rect 10788 13574 10800 13626
rect 10852 13574 10864 13626
rect 10916 13574 17047 13626
rect 17099 13574 17111 13626
rect 17163 13574 17175 13626
rect 17227 13574 17239 13626
rect 17291 13574 17303 13626
rect 17355 13574 23486 13626
rect 23538 13574 23550 13626
rect 23602 13574 23614 13626
rect 23666 13574 23678 13626
rect 23730 13574 23742 13626
rect 23794 13574 26864 13626
rect 1104 13552 26864 13574
rect 3234 13472 3240 13524
rect 3292 13472 3298 13524
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 4154 13472 4160 13524
rect 4212 13472 4218 13524
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 4982 13512 4988 13524
rect 4295 13484 4988 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5534 13472 5540 13524
rect 5592 13472 5598 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 7156 13484 7205 13512
rect 7156 13472 7162 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7193 13475 7251 13481
rect 7558 13472 7564 13524
rect 7616 13472 7622 13524
rect 12345 13515 12403 13521
rect 7944 13484 11928 13512
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 4709 13447 4767 13453
rect 4709 13444 4721 13447
rect 4396 13416 4721 13444
rect 4396 13404 4402 13416
rect 4709 13413 4721 13416
rect 4755 13413 4767 13447
rect 4709 13407 4767 13413
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 4154 13376 4160 13388
rect 3559 13348 4160 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4154 13336 4160 13348
rect 4212 13376 4218 13388
rect 5626 13376 5632 13388
rect 4212 13348 4568 13376
rect 4212 13336 4218 13348
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 1670 13308 1676 13320
rect 1627 13280 1676 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2682 13308 2688 13320
rect 1912 13280 2688 13308
rect 1912 13268 1918 13280
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 4540 13317 4568 13348
rect 5184 13348 5632 13376
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3292 13280 3433 13308
rect 3292 13268 3298 13280
rect 3421 13277 3433 13280
rect 3467 13308 3479 13311
rect 4433 13311 4491 13317
rect 3467 13280 3832 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3804 13249 3832 13280
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 2102 13243 2160 13249
rect 2102 13240 2114 13243
rect 1780 13212 2114 13240
rect 1780 13181 1808 13212
rect 2102 13209 2114 13212
rect 2148 13209 2160 13243
rect 2102 13203 2160 13209
rect 3789 13243 3847 13249
rect 3789 13209 3801 13243
rect 3835 13209 3847 13243
rect 3789 13203 3847 13209
rect 3878 13200 3884 13252
rect 3936 13240 3942 13252
rect 3989 13243 4047 13249
rect 3989 13240 4001 13243
rect 3936 13212 4001 13240
rect 3936 13200 3942 13212
rect 3989 13209 4001 13212
rect 4035 13209 4047 13243
rect 3989 13203 4047 13209
rect 1765 13175 1823 13181
rect 1765 13141 1777 13175
rect 1811 13141 1823 13175
rect 4448 13172 4476 13271
rect 4816 13240 4844 13271
rect 4890 13268 4896 13320
rect 4948 13268 4954 13320
rect 5074 13268 5080 13320
rect 5132 13268 5138 13320
rect 5184 13317 5212 13348
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 7944 13376 7972 13484
rect 8570 13444 8576 13456
rect 8496 13416 8576 13444
rect 7852 13348 7972 13376
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5258 13268 5264 13320
rect 5316 13268 5322 13320
rect 5810 13268 5816 13320
rect 5868 13268 5874 13320
rect 6080 13311 6138 13317
rect 6080 13277 6092 13311
rect 6126 13308 6138 13311
rect 6454 13308 6460 13320
rect 6126 13280 6460 13308
rect 6126 13277 6138 13280
rect 6080 13271 6138 13277
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 7742 13268 7748 13320
rect 7800 13268 7806 13320
rect 7852 13317 7880 13348
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8496 13376 8524 13416
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 8846 13404 8852 13456
rect 8904 13444 8910 13456
rect 8941 13447 8999 13453
rect 8941 13444 8953 13447
rect 8904 13416 8953 13444
rect 8904 13404 8910 13416
rect 8941 13413 8953 13416
rect 8987 13413 8999 13447
rect 11900 13444 11928 13484
rect 12345 13481 12357 13515
rect 12391 13512 12403 13515
rect 12802 13512 12808 13524
rect 12391 13484 12808 13512
rect 12391 13481 12403 13484
rect 12345 13475 12403 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13538 13472 13544 13524
rect 13596 13472 13602 13524
rect 14829 13515 14887 13521
rect 14829 13481 14841 13515
rect 14875 13512 14887 13515
rect 15010 13512 15016 13524
rect 14875 13484 15016 13512
rect 14875 13481 14887 13484
rect 14829 13475 14887 13481
rect 15010 13472 15016 13484
rect 15068 13512 15074 13524
rect 15378 13512 15384 13524
rect 15068 13484 15384 13512
rect 15068 13472 15074 13484
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 18325 13515 18383 13521
rect 18325 13481 18337 13515
rect 18371 13512 18383 13515
rect 18874 13512 18880 13524
rect 18371 13484 18880 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 22094 13512 22100 13524
rect 18984 13484 22100 13512
rect 11900 13416 13216 13444
rect 8941 13407 8999 13413
rect 8168 13348 8524 13376
rect 8168 13336 8174 13348
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 5442 13240 5448 13252
rect 4816 13212 5448 13240
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 7852 13240 7880 13271
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8386 13308 8392 13320
rect 7984 13280 8392 13308
rect 7984 13268 7990 13280
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 8496 13317 8524 13348
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13376 10655 13379
rect 11606 13376 11612 13388
rect 10643 13348 11612 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 11606 13336 11612 13348
rect 11664 13376 11670 13388
rect 12066 13376 12072 13388
rect 11664 13348 12072 13376
rect 11664 13336 11670 13348
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12526 13336 12532 13388
rect 12584 13336 12590 13388
rect 13188 13385 13216 13416
rect 17494 13404 17500 13456
rect 17552 13444 17558 13456
rect 18984 13444 19012 13484
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22649 13515 22707 13521
rect 22649 13481 22661 13515
rect 22695 13512 22707 13515
rect 22830 13512 22836 13524
rect 22695 13484 22836 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 23569 13515 23627 13521
rect 23569 13481 23581 13515
rect 23615 13512 23627 13515
rect 24118 13512 24124 13524
rect 23615 13484 24124 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 23198 13444 23204 13456
rect 17552 13416 19012 13444
rect 22848 13416 23204 13444
rect 17552 13404 17558 13416
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 15749 13379 15807 13385
rect 13219 13348 15056 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 7300 13212 7880 13240
rect 8021 13243 8079 13249
rect 7300 13172 7328 13212
rect 8021 13209 8033 13243
rect 8067 13240 8079 13243
rect 8294 13240 8300 13252
rect 8067 13212 8300 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 8294 13200 8300 13212
rect 8352 13200 8358 13252
rect 4448 13144 7328 13172
rect 1765 13135 1823 13141
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7432 13144 8125 13172
rect 7432 13132 7438 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 8496 13172 8524 13271
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 8846 13308 8852 13320
rect 8803 13280 8852 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 10042 13268 10048 13320
rect 10100 13317 10106 13320
rect 10100 13308 10112 13317
rect 10100 13280 10145 13308
rect 10100 13271 10112 13280
rect 10100 13268 10106 13271
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 13262 13308 13268 13320
rect 12400 13280 13268 13308
rect 12400 13268 12406 13280
rect 13262 13268 13268 13280
rect 13320 13308 13326 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13320 13280 13645 13308
rect 13320 13268 13326 13280
rect 13633 13277 13645 13280
rect 13679 13308 13691 13311
rect 13909 13311 13967 13317
rect 13909 13308 13921 13311
rect 13679 13280 13921 13308
rect 13679 13277 13691 13280
rect 13633 13271 13691 13277
rect 13909 13277 13921 13280
rect 13955 13277 13967 13311
rect 13909 13271 13967 13277
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 14918 13268 14924 13320
rect 14976 13268 14982 13320
rect 15028 13308 15056 13348
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 16114 13376 16120 13388
rect 15795 13348 16120 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 18104 13348 18245 13376
rect 18104 13336 18110 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18598 13336 18604 13388
rect 18656 13336 18662 13388
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 19337 13379 19395 13385
rect 19337 13376 19349 13379
rect 19300 13348 19349 13376
rect 19300 13336 19306 13348
rect 19337 13345 19349 13348
rect 19383 13345 19395 13379
rect 19337 13339 19395 13345
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 20680 13348 21373 13376
rect 20680 13336 20686 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 22848 13320 22876 13416
rect 23198 13404 23204 13416
rect 23256 13404 23262 13456
rect 23842 13404 23848 13456
rect 23900 13404 23906 13456
rect 23934 13404 23940 13456
rect 23992 13404 23998 13456
rect 23014 13336 23020 13388
rect 23072 13376 23078 13388
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 23072 13348 23121 13376
rect 23072 13336 23078 13348
rect 23109 13345 23121 13348
rect 23155 13376 23167 13379
rect 23290 13376 23296 13388
rect 23155 13348 23296 13376
rect 23155 13345 23167 13348
rect 23109 13339 23167 13345
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 23952 13376 23980 13404
rect 23768 13348 23980 13376
rect 18138 13308 18144 13320
rect 15028 13280 18144 13308
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 18690 13268 18696 13320
rect 18748 13268 18754 13320
rect 22830 13268 22836 13320
rect 22888 13268 22894 13320
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13308 23259 13311
rect 23382 13308 23388 13320
rect 23247 13280 23388 13308
rect 23247 13277 23259 13280
rect 23201 13271 23259 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23768 13317 23796 13348
rect 24578 13336 24584 13388
rect 24636 13376 24642 13388
rect 24673 13379 24731 13385
rect 24673 13376 24685 13379
rect 24636 13348 24685 13376
rect 24636 13336 24642 13348
rect 24673 13345 24685 13348
rect 24719 13345 24731 13379
rect 24673 13339 24731 13345
rect 23753 13311 23811 13317
rect 23753 13277 23765 13311
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 24026 13268 24032 13320
rect 24084 13268 24090 13320
rect 10873 13243 10931 13249
rect 10873 13209 10885 13243
rect 10919 13240 10931 13243
rect 11146 13240 11152 13252
rect 10919 13212 11152 13240
rect 10919 13209 10931 13212
rect 10873 13203 10931 13209
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 13817 13243 13875 13249
rect 13817 13240 13829 13243
rect 12098 13212 13829 13240
rect 13817 13209 13829 13212
rect 13863 13209 13875 13243
rect 15746 13240 15752 13252
rect 13817 13203 13875 13209
rect 14936 13212 15752 13240
rect 14936 13172 14964 13212
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 15841 13243 15899 13249
rect 15841 13209 15853 13243
rect 15887 13240 15899 13243
rect 16942 13240 16948 13252
rect 15887 13212 16948 13240
rect 15887 13209 15899 13212
rect 15841 13203 15899 13209
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 19076 13212 19625 13240
rect 8496 13144 14964 13172
rect 8113 13135 8171 13141
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15197 13175 15255 13181
rect 15197 13172 15209 13175
rect 15068 13144 15209 13172
rect 15068 13132 15074 13144
rect 15197 13141 15209 13144
rect 15243 13141 15255 13175
rect 15197 13135 15255 13141
rect 15286 13132 15292 13184
rect 15344 13172 15350 13184
rect 15930 13172 15936 13184
rect 15344 13144 15936 13172
rect 15344 13132 15350 13144
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 16301 13175 16359 13181
rect 16301 13172 16313 13175
rect 16172 13144 16313 13172
rect 16172 13132 16178 13144
rect 16301 13141 16313 13144
rect 16347 13141 16359 13175
rect 16301 13135 16359 13141
rect 17957 13175 18015 13181
rect 17957 13141 17969 13175
rect 18003 13172 18015 13175
rect 18138 13172 18144 13184
rect 18003 13144 18144 13172
rect 18003 13141 18015 13144
rect 17957 13135 18015 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 19076 13181 19104 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 20070 13200 20076 13252
rect 20128 13200 20134 13252
rect 24946 13249 24952 13252
rect 24940 13203 24952 13249
rect 24946 13200 24952 13203
rect 25004 13200 25010 13252
rect 19061 13175 19119 13181
rect 19061 13141 19073 13175
rect 19107 13141 19119 13175
rect 19061 13135 19119 13141
rect 26053 13175 26111 13181
rect 26053 13141 26065 13175
rect 26099 13172 26111 13175
rect 26234 13172 26240 13184
rect 26099 13144 26240 13172
rect 26099 13141 26111 13144
rect 26053 13135 26111 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 1104 13082 26864 13104
rect 1104 13030 4829 13082
rect 4881 13030 4893 13082
rect 4945 13030 4957 13082
rect 5009 13030 5021 13082
rect 5073 13030 5085 13082
rect 5137 13030 11268 13082
rect 11320 13030 11332 13082
rect 11384 13030 11396 13082
rect 11448 13030 11460 13082
rect 11512 13030 11524 13082
rect 11576 13030 17707 13082
rect 17759 13030 17771 13082
rect 17823 13030 17835 13082
rect 17887 13030 17899 13082
rect 17951 13030 17963 13082
rect 18015 13030 24146 13082
rect 24198 13030 24210 13082
rect 24262 13030 24274 13082
rect 24326 13030 24338 13082
rect 24390 13030 24402 13082
rect 24454 13030 26864 13082
rect 1104 13008 26864 13030
rect 3237 12971 3295 12977
rect 3237 12937 3249 12971
rect 3283 12968 3295 12971
rect 3418 12968 3424 12980
rect 3283 12940 3424 12968
rect 3283 12937 3295 12940
rect 3237 12931 3295 12937
rect 3418 12928 3424 12940
rect 3476 12968 3482 12980
rect 3786 12968 3792 12980
rect 3476 12940 3792 12968
rect 3476 12928 3482 12940
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 4893 12971 4951 12977
rect 4893 12968 4905 12971
rect 3936 12940 4905 12968
rect 3936 12928 3942 12940
rect 4893 12937 4905 12940
rect 4939 12937 4951 12971
rect 7558 12968 7564 12980
rect 4893 12931 4951 12937
rect 5184 12940 7564 12968
rect 3970 12860 3976 12912
rect 4028 12860 4034 12912
rect 4338 12860 4344 12912
rect 4396 12900 4402 12912
rect 5184 12900 5212 12940
rect 4396 12872 5212 12900
rect 4396 12860 4402 12872
rect 5258 12860 5264 12912
rect 5316 12860 5322 12912
rect 5368 12909 5396 12940
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 7745 12971 7803 12977
rect 7745 12937 7757 12971
rect 7791 12968 7803 12971
rect 7926 12968 7932 12980
rect 7791 12940 7932 12968
rect 7791 12937 7803 12940
rect 7745 12931 7803 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8021 12971 8079 12977
rect 8021 12937 8033 12971
rect 8067 12968 8079 12971
rect 8570 12968 8576 12980
rect 8067 12940 8576 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 11422 12968 11428 12980
rect 10980 12940 11428 12968
rect 5353 12903 5411 12909
rect 5353 12869 5365 12903
rect 5399 12869 5411 12903
rect 5353 12863 5411 12869
rect 9309 12903 9367 12909
rect 9309 12869 9321 12903
rect 9355 12900 9367 12903
rect 9398 12900 9404 12912
rect 9355 12872 9404 12900
rect 9355 12869 9367 12872
rect 9309 12863 9367 12869
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 10980 12900 11008 12940
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11698 12968 11704 12980
rect 11563 12940 11704 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 12216 12940 12541 12968
rect 12216 12928 12222 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 12529 12931 12587 12937
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 15562 12968 15568 12980
rect 13320 12940 15568 12968
rect 13320 12928 13326 12940
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 17494 12968 17500 12980
rect 15804 12940 17500 12968
rect 15804 12928 15810 12940
rect 17494 12928 17500 12940
rect 17552 12968 17558 12980
rect 17957 12971 18015 12977
rect 17957 12968 17969 12971
rect 17552 12940 17969 12968
rect 17552 12928 17558 12940
rect 17957 12937 17969 12940
rect 18003 12937 18015 12971
rect 17957 12931 18015 12937
rect 19797 12971 19855 12977
rect 19797 12937 19809 12971
rect 19843 12968 19855 12971
rect 20070 12968 20076 12980
rect 19843 12940 20076 12968
rect 19843 12937 19855 12940
rect 19797 12931 19855 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20990 12928 20996 12980
rect 21048 12928 21054 12980
rect 23753 12971 23811 12977
rect 23753 12937 23765 12971
rect 23799 12968 23811 12971
rect 23934 12968 23940 12980
rect 23799 12940 23940 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 24305 12971 24363 12977
rect 24305 12937 24317 12971
rect 24351 12968 24363 12971
rect 24670 12968 24676 12980
rect 24351 12940 24676 12968
rect 24351 12937 24363 12940
rect 24305 12931 24363 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 24857 12971 24915 12977
rect 24857 12937 24869 12971
rect 24903 12968 24915 12971
rect 24946 12968 24952 12980
rect 24903 12940 24952 12968
rect 24903 12937 24915 12940
rect 24857 12931 24915 12937
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 10626 12872 11008 12900
rect 11054 12860 11060 12912
rect 11112 12860 11118 12912
rect 12066 12900 12072 12912
rect 11624 12872 12072 12900
rect 11624 12844 11652 12872
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 13446 12900 13452 12912
rect 12124 12872 13452 12900
rect 12124 12860 12130 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 14737 12903 14795 12909
rect 14737 12869 14749 12903
rect 14783 12900 14795 12903
rect 15470 12900 15476 12912
rect 14783 12872 15476 12900
rect 14783 12869 14795 12872
rect 14737 12863 14795 12869
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 15988 12872 18000 12900
rect 15988 12860 15994 12872
rect 1854 12792 1860 12844
rect 1912 12792 1918 12844
rect 2124 12835 2182 12841
rect 2124 12801 2136 12835
rect 2170 12832 2182 12835
rect 3326 12832 3332 12844
rect 2170 12804 3332 12832
rect 2170 12801 2182 12804
rect 2124 12795 2182 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3418 12792 3424 12844
rect 3476 12792 3482 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4522 12832 4528 12844
rect 4479 12804 4528 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 4632 12764 4660 12792
rect 4540 12736 4660 12764
rect 5184 12764 5212 12795
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5500 12804 5549 12832
rect 5500 12792 5506 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7156 12804 7665 12832
rect 7156 12792 7162 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7892 12804 7941 12832
rect 7892 12792 7898 12804
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 8076 12804 8217 12832
rect 8076 12792 8082 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 8662 12792 8668 12844
rect 8720 12792 8726 12844
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11606 12832 11612 12844
rect 11379 12804 11612 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12250 12832 12256 12844
rect 11931 12804 12256 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13170 12832 13176 12844
rect 12759 12804 13176 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15286 12832 15292 12844
rect 15243 12804 15292 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15580 12804 15669 12832
rect 5626 12764 5632 12776
rect 5184 12736 5632 12764
rect 4540 12705 4568 12736
rect 5626 12724 5632 12736
rect 5684 12764 5690 12776
rect 8110 12764 8116 12776
rect 5684 12736 8116 12764
rect 5684 12724 5690 12736
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 8754 12764 8760 12776
rect 8527 12736 8760 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 9640 12736 11989 12764
rect 9640 12724 9646 12736
rect 11977 12733 11989 12736
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12665 4583 12699
rect 4525 12659 4583 12665
rect 4614 12656 4620 12708
rect 4672 12656 4678 12708
rect 4985 12699 5043 12705
rect 4985 12665 4997 12699
rect 5031 12696 5043 12699
rect 5166 12696 5172 12708
rect 5031 12668 5172 12696
rect 5031 12665 5043 12668
rect 4985 12659 5043 12665
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 8573 12699 8631 12705
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 8619 12668 8861 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 8849 12665 8861 12668
rect 8895 12665 8907 12699
rect 8849 12659 8907 12665
rect 9030 12656 9036 12708
rect 9088 12656 9094 12708
rect 12176 12696 12204 12727
rect 15010 12724 15016 12776
rect 15068 12724 15074 12776
rect 15102 12724 15108 12776
rect 15160 12724 15166 12776
rect 13262 12696 13268 12708
rect 12176 12668 13268 12696
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 15580 12705 15608 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 17972 12832 18000 12872
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 19981 12903 20039 12909
rect 19981 12900 19993 12903
rect 18748 12872 19993 12900
rect 18748 12860 18754 12872
rect 19981 12869 19993 12872
rect 20027 12869 20039 12903
rect 19981 12863 20039 12869
rect 18046 12832 18052 12844
rect 17972 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12832 18110 12844
rect 18877 12835 18935 12841
rect 18877 12832 18889 12835
rect 18104 12804 18889 12832
rect 18104 12792 18110 12804
rect 18877 12801 18889 12804
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12832 19763 12835
rect 20806 12832 20812 12844
rect 19751 12804 20812 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 17865 12767 17923 12773
rect 15672 12736 17816 12764
rect 15565 12699 15623 12705
rect 13372 12668 15516 12696
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4430 12628 4436 12640
rect 4028 12600 4436 12628
rect 4028 12588 4034 12600
rect 4430 12588 4436 12600
rect 4488 12628 4494 12640
rect 9048 12628 9076 12656
rect 4488 12600 9076 12628
rect 4488 12588 4494 12600
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 13372 12628 13400 12668
rect 9180 12600 13400 12628
rect 9180 12588 9186 12600
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 15378 12628 15384 12640
rect 13504 12600 15384 12628
rect 13504 12588 13510 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 15488 12628 15516 12668
rect 15565 12665 15577 12699
rect 15611 12665 15623 12699
rect 15565 12659 15623 12665
rect 15672 12628 15700 12736
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 15933 12699 15991 12705
rect 15933 12696 15945 12699
rect 15804 12668 15945 12696
rect 15804 12656 15810 12668
rect 15933 12665 15945 12668
rect 15979 12665 15991 12699
rect 17788 12696 17816 12736
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18138 12764 18144 12776
rect 17911 12736 18144 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12733 19027 12767
rect 19076 12764 19104 12792
rect 19996 12776 20024 12804
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 19076 12736 19165 12764
rect 18969 12727 19027 12733
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 18984 12696 19012 12727
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 20622 12724 20628 12776
rect 20680 12724 20686 12776
rect 24213 12767 24271 12773
rect 24213 12733 24225 12767
rect 24259 12764 24271 12767
rect 24780 12764 24808 12795
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25038 12832 25044 12844
rect 24912 12804 25044 12832
rect 24912 12792 24918 12804
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25314 12792 25320 12844
rect 25372 12792 25378 12844
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12832 25559 12835
rect 25777 12835 25835 12841
rect 25777 12832 25789 12835
rect 25547 12804 25789 12832
rect 25547 12801 25559 12804
rect 25501 12795 25559 12801
rect 25777 12801 25789 12804
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 26234 12764 26240 12776
rect 24259 12736 26240 12764
rect 24259 12733 24271 12736
rect 24213 12727 24271 12733
rect 26234 12724 26240 12736
rect 26292 12764 26298 12776
rect 26329 12767 26387 12773
rect 26329 12764 26341 12767
rect 26292 12736 26341 12764
rect 26292 12724 26298 12736
rect 26329 12733 26341 12736
rect 26375 12733 26387 12767
rect 26329 12727 26387 12733
rect 20806 12696 20812 12708
rect 17788 12668 20812 12696
rect 15933 12659 15991 12665
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 20990 12656 20996 12708
rect 21048 12696 21054 12708
rect 23845 12699 23903 12705
rect 23845 12696 23857 12699
rect 21048 12668 23857 12696
rect 21048 12656 21054 12668
rect 23845 12665 23857 12668
rect 23891 12696 23903 12699
rect 23891 12668 24532 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 15488 12600 15700 12628
rect 15841 12631 15899 12637
rect 15841 12597 15853 12631
rect 15887 12628 15899 12631
rect 16206 12628 16212 12640
rect 15887 12600 16212 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 18414 12588 18420 12640
rect 18472 12588 18478 12640
rect 18506 12588 18512 12640
rect 18564 12588 18570 12640
rect 21818 12588 21824 12640
rect 21876 12588 21882 12640
rect 24504 12637 24532 12668
rect 24489 12631 24547 12637
rect 24489 12597 24501 12631
rect 24535 12597 24547 12631
rect 24489 12591 24547 12597
rect 1104 12538 26864 12560
rect 1104 12486 4169 12538
rect 4221 12486 4233 12538
rect 4285 12486 4297 12538
rect 4349 12486 4361 12538
rect 4413 12486 4425 12538
rect 4477 12486 10608 12538
rect 10660 12486 10672 12538
rect 10724 12486 10736 12538
rect 10788 12486 10800 12538
rect 10852 12486 10864 12538
rect 10916 12486 17047 12538
rect 17099 12486 17111 12538
rect 17163 12486 17175 12538
rect 17227 12486 17239 12538
rect 17291 12486 17303 12538
rect 17355 12486 23486 12538
rect 23538 12486 23550 12538
rect 23602 12486 23614 12538
rect 23666 12486 23678 12538
rect 23730 12486 23742 12538
rect 23794 12486 26864 12538
rect 1104 12464 26864 12486
rect 3970 12384 3976 12436
rect 4028 12384 4034 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4522 12424 4528 12436
rect 4295 12396 4528 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4672 12396 4721 12424
rect 4672 12384 4678 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 8297 12427 8355 12433
rect 8297 12393 8309 12427
rect 8343 12424 8355 12427
rect 8478 12424 8484 12436
rect 8343 12396 8484 12424
rect 8343 12393 8355 12396
rect 8297 12387 8355 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12802 12424 12808 12436
rect 12391 12396 12808 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 17000 12396 17233 12424
rect 17000 12384 17006 12396
rect 17221 12393 17233 12396
rect 17267 12424 17279 12427
rect 20898 12424 20904 12436
rect 17267 12396 20904 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21634 12384 21640 12436
rect 21692 12424 21698 12436
rect 21913 12427 21971 12433
rect 21692 12396 21864 12424
rect 21692 12384 21698 12396
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 5166 12356 5172 12368
rect 2740 12328 5172 12356
rect 2740 12316 2746 12328
rect 5166 12316 5172 12328
rect 5224 12356 5230 12368
rect 5810 12356 5816 12368
rect 5224 12328 5816 12356
rect 5224 12316 5230 12328
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 8665 12359 8723 12365
rect 8665 12356 8677 12359
rect 8444 12328 8677 12356
rect 8444 12316 8450 12328
rect 8665 12325 8677 12328
rect 8711 12325 8723 12359
rect 8665 12319 8723 12325
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 21729 12359 21787 12365
rect 21729 12356 21741 12359
rect 21416 12328 21741 12356
rect 21416 12316 21422 12328
rect 21729 12325 21741 12328
rect 21775 12325 21787 12359
rect 21836 12356 21864 12396
rect 21913 12393 21925 12427
rect 21959 12424 21971 12427
rect 22002 12424 22008 12436
rect 21959 12396 22008 12424
rect 21959 12393 21971 12396
rect 21913 12387 21971 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22830 12384 22836 12436
rect 22888 12384 22894 12436
rect 22848 12356 22876 12384
rect 23382 12356 23388 12368
rect 21836 12328 23388 12356
rect 21729 12319 21787 12325
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3418 12288 3424 12300
rect 2915 12260 3424 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 4212 12260 4353 12288
rect 4212 12248 4218 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 8205 12291 8263 12297
rect 8205 12288 8217 12291
rect 7432 12260 8217 12288
rect 7432 12248 7438 12260
rect 8205 12257 8217 12260
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15436 12260 15485 12288
rect 15436 12248 15442 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15746 12248 15752 12300
rect 15804 12248 15810 12300
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 17644 12260 18153 12288
rect 17644 12248 17650 12260
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 19058 12248 19064 12300
rect 19116 12288 19122 12300
rect 19116 12260 20760 12288
rect 19116 12248 19122 12260
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2133 12223 2191 12229
rect 2133 12220 2145 12223
rect 2096 12192 2145 12220
rect 2096 12180 2102 12192
rect 2133 12189 2145 12192
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2314 12220 2320 12232
rect 2271 12192 2320 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2455 12192 2774 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2746 12152 2774 12192
rect 3786 12180 3792 12232
rect 3844 12180 3850 12232
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 7650 12220 7656 12232
rect 4571 12192 7656 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8352 12192 8493 12220
rect 8352 12180 8358 12192
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11790 12220 11796 12232
rect 11563 12192 11796 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11790 12180 11796 12192
rect 11848 12220 11854 12232
rect 12342 12220 12348 12232
rect 11848 12192 12348 12220
rect 11848 12180 11854 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14642 12220 14648 12232
rect 13771 12192 14648 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18046 12220 18052 12232
rect 18003 12192 18052 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 18840 12192 18889 12220
rect 18840 12180 18846 12192
rect 18877 12189 18889 12192
rect 18923 12220 18935 12223
rect 18923 12192 19196 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 9582 12152 9588 12164
rect 2746 12124 9588 12152
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 13480 12155 13538 12161
rect 13480 12121 13492 12155
rect 13526 12121 13538 12155
rect 13480 12115 13538 12121
rect 13495 12084 13523 12115
rect 16758 12112 16764 12164
rect 16816 12112 16822 12164
rect 19058 12152 19064 12164
rect 17236 12124 19064 12152
rect 17236 12084 17264 12124
rect 19058 12112 19064 12124
rect 19116 12112 19122 12164
rect 19168 12152 19196 12192
rect 19242 12180 19248 12232
rect 19300 12180 19306 12232
rect 20732 12220 20760 12260
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 21269 12291 21327 12297
rect 21269 12288 21281 12291
rect 20864 12260 21281 12288
rect 20864 12248 20870 12260
rect 21269 12257 21281 12260
rect 21315 12288 21327 12291
rect 23014 12288 23020 12300
rect 21315 12260 23020 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 21818 12220 21824 12232
rect 20732 12192 21824 12220
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 23106 12180 23112 12232
rect 23164 12180 23170 12232
rect 19426 12152 19432 12164
rect 19168 12124 19432 12152
rect 19426 12112 19432 12124
rect 19484 12112 19490 12164
rect 19518 12112 19524 12164
rect 19576 12112 19582 12164
rect 20070 12112 20076 12164
rect 20128 12112 20134 12164
rect 21450 12112 21456 12164
rect 21508 12112 21514 12164
rect 13495 12056 17264 12084
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17368 12056 17601 12084
rect 17368 12044 17374 12056
rect 17589 12053 17601 12056
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18230 12084 18236 12096
rect 18104 12056 18236 12084
rect 18104 12044 18110 12056
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 18874 12084 18880 12096
rect 18831 12056 18880 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 22646 12044 22652 12096
rect 22704 12044 22710 12096
rect 1104 11994 26864 12016
rect 1104 11942 4829 11994
rect 4881 11942 4893 11994
rect 4945 11942 4957 11994
rect 5009 11942 5021 11994
rect 5073 11942 5085 11994
rect 5137 11942 11268 11994
rect 11320 11942 11332 11994
rect 11384 11942 11396 11994
rect 11448 11942 11460 11994
rect 11512 11942 11524 11994
rect 11576 11942 17707 11994
rect 17759 11942 17771 11994
rect 17823 11942 17835 11994
rect 17887 11942 17899 11994
rect 17951 11942 17963 11994
rect 18015 11942 24146 11994
rect 24198 11942 24210 11994
rect 24262 11942 24274 11994
rect 24326 11942 24338 11994
rect 24390 11942 24402 11994
rect 24454 11942 26864 11994
rect 1104 11920 26864 11942
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14458 11880 14464 11892
rect 14047 11852 14464 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14458 11840 14464 11852
rect 14516 11880 14522 11892
rect 15286 11880 15292 11892
rect 14516 11852 15292 11880
rect 14516 11840 14522 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 16758 11840 16764 11892
rect 16816 11840 16822 11892
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11849 17555 11883
rect 17497 11843 17555 11849
rect 15930 11812 15936 11824
rect 15778 11784 15936 11812
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 16114 11772 16120 11824
rect 16172 11812 16178 11824
rect 16209 11815 16267 11821
rect 16209 11812 16221 11815
rect 16172 11784 16221 11812
rect 16172 11772 16178 11784
rect 16209 11781 16221 11784
rect 16255 11781 16267 11815
rect 17512 11812 17540 11843
rect 18046 11840 18052 11892
rect 18104 11880 18110 11892
rect 18104 11852 19656 11880
rect 18104 11840 18110 11852
rect 17865 11815 17923 11821
rect 17865 11812 17877 11815
rect 17512 11784 17877 11812
rect 16209 11775 16267 11781
rect 17865 11781 17877 11784
rect 17911 11781 17923 11815
rect 17865 11775 17923 11781
rect 18874 11772 18880 11824
rect 18932 11772 18938 11824
rect 19628 11821 19656 11852
rect 20070 11840 20076 11892
rect 20128 11840 20134 11892
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 20956 11852 23888 11880
rect 20956 11840 20962 11852
rect 19613 11815 19671 11821
rect 19613 11781 19625 11815
rect 19659 11812 19671 11815
rect 21634 11812 21640 11824
rect 19659 11784 21640 11812
rect 19659 11781 19671 11784
rect 19613 11775 19671 11781
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 21726 11772 21732 11824
rect 21784 11812 21790 11824
rect 22370 11812 22376 11824
rect 21784 11784 22376 11812
rect 21784 11772 21790 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13219 11716 13676 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13648 11617 13676 11716
rect 16850 11704 16856 11756
rect 16908 11704 16914 11756
rect 17310 11704 17316 11756
rect 17368 11704 17374 11756
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 19978 11744 19984 11756
rect 19484 11716 19984 11744
rect 19484 11704 19490 11716
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11744 21971 11747
rect 22002 11744 22008 11756
rect 21959 11716 22008 11744
rect 21959 11713 21971 11716
rect 21913 11707 21971 11713
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22112 11753 22140 11784
rect 22370 11772 22376 11784
rect 22428 11772 22434 11824
rect 22557 11815 22615 11821
rect 22557 11781 22569 11815
rect 22603 11812 22615 11815
rect 22603 11784 22876 11812
rect 22603 11781 22615 11784
rect 22557 11775 22615 11781
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22462 11744 22468 11756
rect 22327 11716 22468 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 22646 11704 22652 11756
rect 22704 11704 22710 11756
rect 22848 11753 22876 11784
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 23014 11704 23020 11756
rect 23072 11704 23078 11756
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11744 23443 11747
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23431 11716 23673 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 13780 11648 14105 11676
rect 13780 11636 13786 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 14461 11679 14519 11685
rect 14323 11648 14412 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 13633 11611 13691 11617
rect 13633 11577 13645 11611
rect 13679 11577 13691 11611
rect 13633 11571 13691 11577
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12989 11543 13047 11549
rect 12989 11540 13001 11543
rect 12400 11512 13001 11540
rect 12400 11500 12406 11512
rect 12989 11509 13001 11512
rect 13035 11509 13047 11543
rect 14384 11540 14412 11648
rect 14461 11645 14473 11679
rect 14507 11676 14519 11679
rect 14550 11676 14556 11688
rect 14507 11648 14556 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 14550 11636 14556 11648
rect 14608 11676 14614 11688
rect 14608 11648 16436 11676
rect 14608 11636 14614 11648
rect 16408 11608 16436 11648
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 16540 11648 17601 11676
rect 16540 11636 16546 11648
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 22922 11636 22928 11688
rect 22980 11636 22986 11688
rect 23860 11676 23888 11852
rect 24673 11815 24731 11821
rect 24673 11781 24685 11815
rect 24719 11812 24731 11815
rect 24719 11784 25268 11812
rect 24719 11781 24731 11784
rect 24673 11775 24731 11781
rect 25240 11753 25268 11784
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11744 23995 11747
rect 25225 11747 25283 11753
rect 23983 11716 24808 11744
rect 23983 11713 23995 11716
rect 23937 11707 23995 11713
rect 24780 11685 24808 11716
rect 25225 11713 25237 11747
rect 25271 11744 25283 11747
rect 25774 11744 25780 11756
rect 25271 11716 25780 11744
rect 25271 11713 25283 11716
rect 25225 11707 25283 11713
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 26510 11704 26516 11756
rect 26568 11704 26574 11756
rect 24765 11679 24823 11685
rect 23860 11648 24348 11676
rect 16408 11580 16804 11608
rect 16666 11540 16672 11552
rect 14384 11512 16672 11540
rect 12989 11503 13047 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16776 11540 16804 11580
rect 21450 11568 21456 11620
rect 21508 11608 21514 11620
rect 21818 11608 21824 11620
rect 21508 11580 21824 11608
rect 21508 11568 21514 11580
rect 21818 11568 21824 11580
rect 21876 11608 21882 11620
rect 24320 11617 24348 11648
rect 24765 11645 24777 11679
rect 24811 11645 24823 11679
rect 24765 11639 24823 11645
rect 23477 11611 23535 11617
rect 23477 11608 23489 11611
rect 21876 11580 23489 11608
rect 21876 11568 21882 11580
rect 23477 11577 23489 11580
rect 23523 11577 23535 11611
rect 23477 11571 23535 11577
rect 23753 11611 23811 11617
rect 23753 11577 23765 11611
rect 23799 11577 23811 11611
rect 23753 11571 23811 11577
rect 23845 11611 23903 11617
rect 23845 11577 23857 11611
rect 23891 11608 23903 11611
rect 24213 11611 24271 11617
rect 24213 11608 24225 11611
rect 23891 11580 24225 11608
rect 23891 11577 23903 11580
rect 23845 11571 23903 11577
rect 24213 11577 24225 11580
rect 24259 11577 24271 11611
rect 24213 11571 24271 11577
rect 24305 11611 24363 11617
rect 24305 11577 24317 11611
rect 24351 11608 24363 11611
rect 24351 11580 24992 11608
rect 24351 11577 24363 11580
rect 24305 11571 24363 11577
rect 21726 11540 21732 11552
rect 16776 11512 21732 11540
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 23768 11540 23796 11571
rect 23934 11540 23940 11552
rect 23768 11512 23940 11540
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 24964 11549 24992 11580
rect 24949 11543 25007 11549
rect 24949 11509 24961 11543
rect 24995 11509 25007 11543
rect 24949 11503 25007 11509
rect 26326 11500 26332 11552
rect 26384 11500 26390 11552
rect 1104 11450 26864 11472
rect 1104 11398 4169 11450
rect 4221 11398 4233 11450
rect 4285 11398 4297 11450
rect 4349 11398 4361 11450
rect 4413 11398 4425 11450
rect 4477 11398 10608 11450
rect 10660 11398 10672 11450
rect 10724 11398 10736 11450
rect 10788 11398 10800 11450
rect 10852 11398 10864 11450
rect 10916 11398 17047 11450
rect 17099 11398 17111 11450
rect 17163 11398 17175 11450
rect 17227 11398 17239 11450
rect 17291 11398 17303 11450
rect 17355 11398 23486 11450
rect 23538 11398 23550 11450
rect 23602 11398 23614 11450
rect 23666 11398 23678 11450
rect 23730 11398 23742 11450
rect 23794 11398 26864 11450
rect 1104 11376 26864 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 9214 11336 9220 11348
rect 1627 11308 9220 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 11532 11308 15884 11336
rect 3510 11228 3516 11280
rect 3568 11228 3574 11280
rect 3528 11200 3556 11228
rect 4062 11200 4068 11212
rect 3252 11172 4068 11200
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 3252 11141 3280 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5442 11200 5448 11212
rect 5224 11172 5448 11200
rect 5224 11160 5230 11172
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 8570 11200 8576 11212
rect 6963 11172 8576 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 11146 11132 11152 11144
rect 10183 11104 11152 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 3528 11064 3556 11095
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11532 11141 11560 11308
rect 15856 11268 15884 11308
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 15988 11308 16129 11336
rect 15988 11296 15994 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 19518 11336 19524 11348
rect 18739 11308 19524 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 22002 11296 22008 11348
rect 22060 11296 22066 11348
rect 22186 11296 22192 11348
rect 22244 11336 22250 11348
rect 22738 11336 22744 11348
rect 22244 11308 22744 11336
rect 22244 11296 22250 11308
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 22922 11296 22928 11348
rect 22980 11296 22986 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23661 11339 23719 11345
rect 23256 11308 23612 11336
rect 23256 11296 23262 11308
rect 16022 11268 16028 11280
rect 15856 11240 16028 11268
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 18325 11271 18383 11277
rect 18325 11237 18337 11271
rect 18371 11268 18383 11271
rect 18371 11240 19380 11268
rect 18371 11237 18383 11240
rect 18325 11231 18383 11237
rect 11790 11160 11796 11212
rect 11848 11160 11854 11212
rect 12066 11160 12072 11212
rect 12124 11160 12130 11212
rect 12342 11160 12348 11212
rect 12400 11160 12406 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15620 11172 15945 11200
rect 15620 11160 15626 11172
rect 15933 11169 15945 11172
rect 15979 11200 15991 11203
rect 16482 11200 16488 11212
rect 15979 11172 16488 11200
rect 15979 11169 15991 11172
rect 15933 11163 15991 11169
rect 16482 11160 16488 11172
rect 16540 11200 16546 11212
rect 19242 11200 19248 11212
rect 16540 11172 19248 11200
rect 16540 11160 16546 11172
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 19352 11200 19380 11240
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19352 11172 19533 11200
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 21269 11203 21327 11209
rect 21269 11169 21281 11203
rect 21315 11200 21327 11203
rect 22186 11200 22192 11212
rect 21315 11172 22192 11200
rect 21315 11169 21327 11172
rect 21269 11163 21327 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 23216 11200 23244 11296
rect 23382 11228 23388 11280
rect 23440 11268 23446 11280
rect 23477 11271 23535 11277
rect 23477 11268 23489 11271
rect 23440 11240 23489 11268
rect 23440 11228 23446 11240
rect 23477 11237 23489 11240
rect 23523 11237 23535 11271
rect 23584 11268 23612 11308
rect 23661 11305 23673 11339
rect 23707 11336 23719 11339
rect 23934 11336 23940 11348
rect 23707 11308 23940 11336
rect 23707 11305 23719 11308
rect 23661 11299 23719 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 23845 11271 23903 11277
rect 23845 11268 23857 11271
rect 23584 11240 23857 11268
rect 23477 11231 23535 11237
rect 23845 11237 23857 11240
rect 23891 11237 23903 11271
rect 23845 11231 23903 11237
rect 22388 11172 23244 11200
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 3878 11064 3884 11076
rect 3016 11036 3884 11064
rect 3016 11024 3022 11036
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 5408 11036 5457 11064
rect 5408 11024 5414 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 6454 11024 6460 11076
rect 6512 11024 6518 11076
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11532 11064 11560 11095
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 18414 11132 18420 11144
rect 18187 11104 18420 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22388 11141 22416 11172
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 22649 11135 22707 11141
rect 22649 11132 22661 11135
rect 22520 11104 22661 11132
rect 22520 11092 22526 11104
rect 22649 11101 22661 11104
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11132 23995 11135
rect 24578 11132 24584 11144
rect 23983 11104 24584 11132
rect 23983 11101 23995 11104
rect 23937 11095 23995 11101
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 25501 11135 25559 11141
rect 25501 11101 25513 11135
rect 25547 11132 25559 11135
rect 25774 11132 25780 11144
rect 25547 11104 25780 11132
rect 25547 11101 25559 11104
rect 25501 11095 25559 11101
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 11112 11036 11560 11064
rect 11112 11024 11118 11036
rect 13078 11024 13084 11076
rect 13136 11024 13142 11076
rect 15654 11024 15660 11076
rect 15712 11024 15718 11076
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 22557 11067 22615 11073
rect 19668 11036 20010 11064
rect 19668 11024 19674 11036
rect 22557 11033 22569 11067
rect 22603 11064 22615 11067
rect 23014 11064 23020 11076
rect 22603 11036 23020 11064
rect 22603 11033 22615 11036
rect 22557 11027 22615 11033
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 23198 11024 23204 11076
rect 23256 11024 23262 11076
rect 3418 10956 3424 11008
rect 3476 10956 3482 11008
rect 3896 10996 3924 11024
rect 6362 10996 6368 11008
rect 3896 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 8754 10996 8760 11008
rect 6788 10968 8760 10996
rect 6788 10956 6794 10968
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10045 10999 10103 11005
rect 10045 10996 10057 10999
rect 10008 10968 10057 10996
rect 10008 10956 10014 10968
rect 10045 10965 10057 10968
rect 10091 10965 10103 10999
rect 10045 10959 10103 10965
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 13817 10999 13875 11005
rect 13817 10996 13829 10999
rect 13688 10968 13829 10996
rect 13688 10956 13694 10968
rect 13817 10965 13829 10968
rect 13863 10965 13875 10999
rect 13817 10959 13875 10965
rect 14182 10956 14188 11008
rect 14240 10956 14246 11008
rect 24854 10956 24860 11008
rect 24912 10956 24918 11008
rect 1104 10906 26864 10928
rect 1104 10854 4829 10906
rect 4881 10854 4893 10906
rect 4945 10854 4957 10906
rect 5009 10854 5021 10906
rect 5073 10854 5085 10906
rect 5137 10854 11268 10906
rect 11320 10854 11332 10906
rect 11384 10854 11396 10906
rect 11448 10854 11460 10906
rect 11512 10854 11524 10906
rect 11576 10854 17707 10906
rect 17759 10854 17771 10906
rect 17823 10854 17835 10906
rect 17887 10854 17899 10906
rect 17951 10854 17963 10906
rect 18015 10854 24146 10906
rect 24198 10854 24210 10906
rect 24262 10854 24274 10906
rect 24326 10854 24338 10906
rect 24390 10854 24402 10906
rect 24454 10854 26864 10906
rect 1104 10832 26864 10854
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 5258 10792 5264 10804
rect 4304 10764 5264 10792
rect 4304 10752 4310 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 8018 10792 8024 10804
rect 6564 10764 8024 10792
rect 1854 10724 1860 10736
rect 1596 10696 1860 10724
rect 1596 10665 1624 10696
rect 1854 10684 1860 10696
rect 1912 10684 1918 10736
rect 3418 10724 3424 10736
rect 3082 10696 3424 10724
rect 3418 10684 3424 10696
rect 3476 10684 3482 10736
rect 5534 10724 5540 10736
rect 3528 10696 5540 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 3528 10588 3556 10696
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 3878 10616 3884 10668
rect 3936 10616 3942 10668
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 4028 10628 4077 10656
rect 4028 10616 4034 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4387 10628 4813 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4801 10625 4813 10628
rect 4847 10656 4859 10659
rect 4890 10656 4896 10668
rect 4847 10628 4896 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5258 10656 5264 10668
rect 5123 10628 5264 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 1903 10560 3556 10588
rect 3605 10591 3663 10597
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 4264 10588 4292 10616
rect 3651 10560 4292 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5000 10588 5028 10619
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5902 10656 5908 10668
rect 5675 10628 5908 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 4672 10560 5028 10588
rect 5368 10588 5396 10619
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 6564 10665 6592 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8662 10792 8668 10804
rect 8168 10764 8668 10792
rect 8168 10752 8174 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8812 10764 10640 10792
rect 8812 10752 8818 10764
rect 6822 10684 6828 10736
rect 6880 10724 6886 10736
rect 7561 10727 7619 10733
rect 7561 10724 7573 10727
rect 6880 10696 7573 10724
rect 6880 10684 6886 10696
rect 7561 10693 7573 10696
rect 7607 10693 7619 10727
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 7561 10687 7619 10693
rect 7668 10696 8401 10724
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6420 10628 6561 10656
rect 6420 10616 6426 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 7668 10656 7696 10696
rect 8389 10693 8401 10696
rect 8435 10724 8447 10727
rect 9398 10724 9404 10736
rect 8435 10696 9404 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 9398 10684 9404 10696
rect 9456 10684 9462 10736
rect 10612 10724 10640 10764
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11204 10764 11529 10792
rect 11204 10752 11210 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 13078 10752 13084 10804
rect 13136 10792 13142 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 13136 10764 13185 10792
rect 13136 10752 13142 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 15654 10792 15660 10804
rect 14047 10764 15660 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 19610 10752 19616 10804
rect 19668 10752 19674 10804
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 22612 10764 22845 10792
rect 22612 10752 22618 10764
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 24854 10792 24860 10804
rect 22833 10755 22891 10761
rect 23860 10764 24860 10792
rect 10612 10696 14320 10724
rect 7524 10628 7696 10656
rect 7524 10616 7530 10628
rect 8110 10616 8116 10668
rect 8168 10616 8174 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8570 10656 8576 10668
rect 8527 10628 8576 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8662 10616 8668 10668
rect 8720 10616 8726 10668
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 11204 10628 11345 10656
rect 11204 10616 11210 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 11848 10628 13093 10656
rect 11848 10616 11854 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14292 10656 14320 10696
rect 14458 10684 14464 10736
rect 14516 10724 14522 10736
rect 14553 10727 14611 10733
rect 14553 10724 14565 10727
rect 14516 10696 14565 10724
rect 14516 10684 14522 10696
rect 14553 10693 14565 10696
rect 14599 10693 14611 10727
rect 14553 10687 14611 10693
rect 21818 10684 21824 10736
rect 21876 10724 21882 10736
rect 22433 10727 22491 10733
rect 22433 10724 22445 10727
rect 21876 10696 22445 10724
rect 21876 10684 21882 10696
rect 22433 10693 22445 10696
rect 22479 10693 22491 10727
rect 22433 10687 22491 10693
rect 22649 10727 22707 10733
rect 22649 10693 22661 10727
rect 22695 10693 22707 10727
rect 22649 10687 22707 10693
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 13863 10628 14228 10656
rect 14292 10628 15025 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 5368 10560 5672 10588
rect 4672 10548 4678 10560
rect 5644 10532 5672 10560
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 6972 10560 8309 10588
rect 6972 10548 6978 10560
rect 8297 10557 8309 10560
rect 8343 10588 8355 10591
rect 8938 10588 8944 10600
rect 8343 10560 8944 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9030 10548 9036 10600
rect 9088 10548 9094 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 9140 10560 9321 10588
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 4157 10523 4215 10529
rect 4157 10520 4169 10523
rect 4120 10492 4169 10520
rect 4120 10480 4126 10492
rect 4157 10489 4169 10492
rect 4203 10489 4215 10523
rect 4157 10483 4215 10489
rect 4525 10523 4583 10529
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 4706 10520 4712 10532
rect 4571 10492 4712 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 5132 10492 5304 10520
rect 5132 10480 5138 10492
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3752 10424 3801 10452
rect 3752 10412 3758 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 4614 10412 4620 10464
rect 4672 10412 4678 10464
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 5276 10452 5304 10492
rect 5350 10480 5356 10532
rect 5408 10480 5414 10532
rect 5626 10480 5632 10532
rect 5684 10480 5690 10532
rect 7929 10523 7987 10529
rect 7929 10520 7941 10523
rect 5980 10492 7941 10520
rect 5980 10452 6008 10492
rect 7929 10489 7941 10492
rect 7975 10520 7987 10523
rect 8202 10520 8208 10532
rect 7975 10492 8208 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 8570 10520 8576 10532
rect 8404 10492 8576 10520
rect 5276 10424 6008 10452
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 7834 10452 7840 10464
rect 7791 10424 7840 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8404 10461 8432 10492
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 9140 10520 9168 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 9456 10560 11069 10588
rect 9456 10548 9462 10560
rect 11057 10557 11069 10560
rect 11103 10588 11115 10591
rect 11698 10588 11704 10600
rect 11103 10560 11704 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12066 10548 12072 10600
rect 12124 10548 12130 10600
rect 14200 10529 14228 10628
rect 15013 10625 15025 10628
rect 15059 10656 15071 10659
rect 15286 10656 15292 10668
rect 15059 10628 15292 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 19484 10628 19533 10656
rect 19484 10616 19490 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22094 10656 22100 10668
rect 22051 10628 22100 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22094 10616 22100 10628
rect 22152 10656 22158 10668
rect 22664 10656 22692 10687
rect 22922 10656 22928 10668
rect 22152 10628 22508 10656
rect 22664 10628 22928 10656
rect 22152 10616 22158 10628
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14516 10560 14657 10588
rect 14516 10548 14522 10560
rect 14645 10557 14657 10560
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 14734 10548 14740 10600
rect 14792 10548 14798 10600
rect 15194 10548 15200 10600
rect 15252 10548 15258 10600
rect 8812 10492 9168 10520
rect 14185 10523 14243 10529
rect 8812 10480 8818 10492
rect 14185 10489 14197 10523
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10421 8447 10455
rect 8389 10415 8447 10421
rect 8478 10412 8484 10464
rect 8536 10412 8542 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9490 10452 9496 10464
rect 8720 10424 9496 10452
rect 8720 10412 8726 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 22186 10412 22192 10464
rect 22244 10412 22250 10464
rect 22278 10412 22284 10464
rect 22336 10412 22342 10464
rect 22480 10461 22508 10628
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 23860 10665 23888 10764
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 25774 10752 25780 10804
rect 25832 10752 25838 10804
rect 24305 10727 24363 10733
rect 24305 10693 24317 10727
rect 24351 10724 24363 10727
rect 24642 10727 24700 10733
rect 24642 10724 24654 10727
rect 24351 10696 24654 10724
rect 24351 10693 24363 10696
rect 24305 10687 24363 10693
rect 24642 10693 24654 10696
rect 24688 10693 24700 10727
rect 24642 10687 24700 10693
rect 23845 10659 23903 10665
rect 23845 10625 23857 10659
rect 23891 10625 23903 10659
rect 23845 10619 23903 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10656 24455 10659
rect 24486 10656 24492 10668
rect 24443 10628 24492 10656
rect 24443 10625 24455 10628
rect 24397 10619 24455 10625
rect 22465 10455 22523 10461
rect 22465 10421 22477 10455
rect 22511 10452 22523 10455
rect 22738 10452 22744 10464
rect 22511 10424 22744 10452
rect 22511 10421 22523 10424
rect 22465 10415 22523 10421
rect 22738 10412 22744 10424
rect 22796 10412 22802 10464
rect 23937 10455 23995 10461
rect 23937 10421 23949 10455
rect 23983 10452 23995 10455
rect 24026 10452 24032 10464
rect 23983 10424 24032 10452
rect 23983 10421 23995 10424
rect 23937 10415 23995 10421
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24136 10452 24164 10619
rect 24486 10616 24492 10628
rect 24544 10616 24550 10668
rect 25038 10452 25044 10464
rect 24136 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 1104 10362 26864 10384
rect 1104 10310 4169 10362
rect 4221 10310 4233 10362
rect 4285 10310 4297 10362
rect 4349 10310 4361 10362
rect 4413 10310 4425 10362
rect 4477 10310 10608 10362
rect 10660 10310 10672 10362
rect 10724 10310 10736 10362
rect 10788 10310 10800 10362
rect 10852 10310 10864 10362
rect 10916 10310 17047 10362
rect 17099 10310 17111 10362
rect 17163 10310 17175 10362
rect 17227 10310 17239 10362
rect 17291 10310 17303 10362
rect 17355 10310 23486 10362
rect 23538 10310 23550 10362
rect 23602 10310 23614 10362
rect 23666 10310 23678 10362
rect 23730 10310 23742 10362
rect 23794 10310 26864 10362
rect 1104 10288 26864 10310
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 5074 10248 5080 10260
rect 4120 10220 5080 10248
rect 4120 10208 4126 10220
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 5626 10208 5632 10260
rect 5684 10208 5690 10260
rect 7742 10248 7748 10260
rect 5736 10220 7748 10248
rect 4614 10140 4620 10192
rect 4672 10140 4678 10192
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1854 10112 1860 10124
rect 1627 10084 1860 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 4632 10112 4660 10140
rect 4172 10084 4660 10112
rect 4172 10053 4200 10084
rect 5074 10072 5080 10124
rect 5132 10072 5138 10124
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 5736 10112 5764 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8297 10251 8355 10257
rect 8297 10217 8309 10251
rect 8343 10248 8355 10251
rect 8754 10248 8760 10260
rect 8343 10220 8760 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 9548 10220 11437 10248
rect 9548 10208 9554 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 12066 10248 12072 10260
rect 11471 10220 12072 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 14550 10208 14556 10260
rect 14608 10208 14614 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 21876 10220 22140 10248
rect 21876 10208 21882 10220
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6822 10180 6828 10192
rect 5868 10152 6828 10180
rect 5868 10140 5874 10152
rect 6822 10140 6828 10152
rect 6880 10140 6886 10192
rect 8478 10180 8484 10192
rect 7392 10152 8484 10180
rect 7392 10121 7420 10152
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 9263 10183 9321 10189
rect 9263 10180 9275 10183
rect 8628 10152 9275 10180
rect 8628 10140 8634 10152
rect 9263 10149 9275 10152
rect 9309 10149 9321 10183
rect 9263 10143 9321 10149
rect 13722 10140 13728 10192
rect 13780 10140 13786 10192
rect 14369 10183 14427 10189
rect 14369 10149 14381 10183
rect 14415 10180 14427 10183
rect 14458 10180 14464 10192
rect 14415 10152 14464 10180
rect 14415 10149 14427 10152
rect 14369 10143 14427 10149
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 22005 10183 22063 10189
rect 22005 10149 22017 10183
rect 22051 10149 22063 10183
rect 22112 10180 22140 10220
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22244 10220 22293 10248
rect 22244 10208 22250 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 22370 10208 22376 10260
rect 22428 10248 22434 10260
rect 22428 10220 24440 10248
rect 22428 10208 22434 10220
rect 22112 10152 22968 10180
rect 22005 10143 22063 10149
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 5316 10084 5764 10112
rect 5316 10072 5322 10084
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4856 10016 4905 10044
rect 4856 10004 4862 10016
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 5166 10004 5172 10056
rect 5224 10004 5230 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9945 1915 9979
rect 1857 9939 1915 9945
rect 1872 9908 1900 9939
rect 2866 9936 2872 9988
rect 2924 9936 2930 9988
rect 3605 9979 3663 9985
rect 3605 9945 3617 9979
rect 3651 9976 3663 9979
rect 3651 9948 4200 9976
rect 3651 9945 3663 9948
rect 3605 9939 3663 9945
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 1872 9880 3985 9908
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 4172 9908 4200 9948
rect 4246 9936 4252 9988
rect 4304 9936 4310 9988
rect 4338 9936 4344 9988
rect 4396 9936 4402 9988
rect 4479 9979 4537 9985
rect 4479 9945 4491 9979
rect 4525 9976 4537 9979
rect 4709 9979 4767 9985
rect 4709 9976 4721 9979
rect 4525 9948 4721 9976
rect 4525 9945 4537 9948
rect 4479 9939 4537 9945
rect 4709 9945 4721 9948
rect 4755 9976 4767 9979
rect 5368 9976 5396 10007
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 5736 10044 5764 10084
rect 6288 10084 7389 10112
rect 5675 10016 5764 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 6288 10053 6316 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 7699 10084 8156 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5960 10016 6101 10044
rect 5960 10004 5966 10016
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 5813 9979 5871 9985
rect 5813 9976 5825 9979
rect 4755 9948 5825 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 5813 9945 5825 9948
rect 5859 9976 5871 9979
rect 6362 9976 6368 9988
rect 5859 9948 6368 9976
rect 5859 9945 5871 9948
rect 5813 9939 5871 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 6454 9936 6460 9988
rect 6512 9936 6518 9988
rect 6564 9976 6592 10007
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7466 10044 7472 10056
rect 7331 10016 7472 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 8128 10053 8156 10084
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9088 10084 9689 10112
rect 9088 10072 9094 10084
rect 9677 10081 9689 10084
rect 9723 10112 9735 10115
rect 10318 10112 10324 10124
rect 9723 10084 10324 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10318 10072 10324 10084
rect 10376 10112 10382 10124
rect 11609 10115 11667 10121
rect 11609 10112 11621 10115
rect 10376 10084 11621 10112
rect 10376 10072 10382 10084
rect 11609 10081 11621 10084
rect 11655 10081 11667 10115
rect 22020 10112 22048 10143
rect 22738 10112 22744 10124
rect 22020 10084 22744 10112
rect 11609 10075 11667 10081
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7892 10016 7941 10044
rect 7892 10004 7898 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8260 10016 8401 10044
rect 8260 10004 8266 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 7558 9976 7564 9988
rect 6564 9948 7564 9976
rect 7558 9936 7564 9948
rect 7616 9936 7622 9988
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9945 8079 9979
rect 8588 9976 8616 10007
rect 8938 10004 8944 10056
rect 8996 10004 9002 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9306 10044 9312 10056
rect 9171 10016 9312 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9490 10044 9496 10056
rect 9447 10016 9496 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 13630 10044 13636 10056
rect 13587 10016 13636 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14182 10004 14188 10056
rect 14240 10004 14246 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 15194 10044 15200 10056
rect 14507 10016 15200 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 22940 10053 22968 10152
rect 24412 10053 24440 10220
rect 24486 10072 24492 10124
rect 24544 10112 24550 10124
rect 24673 10115 24731 10121
rect 24673 10112 24685 10115
rect 24544 10084 24685 10112
rect 24544 10072 24550 10084
rect 24673 10081 24685 10084
rect 24719 10081 24731 10115
rect 24673 10075 24731 10081
rect 20625 10047 20683 10053
rect 20625 10044 20637 10047
rect 19484 10016 20637 10044
rect 19484 10004 19490 10016
rect 20625 10013 20637 10016
rect 20671 10013 20683 10047
rect 20625 10007 20683 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 8588 9948 9045 9976
rect 8021 9939 8079 9945
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 9033 9939 9091 9945
rect 4982 9908 4988 9920
rect 4172 9880 4988 9908
rect 3973 9871 4031 9877
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6052 9880 6653 9908
rect 6052 9868 6058 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 6641 9871 6699 9877
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9908 7067 9911
rect 7834 9908 7840 9920
rect 7055 9880 7840 9908
rect 7055 9877 7067 9880
rect 7009 9871 7067 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8036 9908 8064 9939
rect 9950 9936 9956 9988
rect 10008 9936 10014 9988
rect 11238 9976 11244 9988
rect 11178 9948 11244 9976
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 11348 9948 11560 9976
rect 7984 9880 8064 9908
rect 7984 9868 7990 9880
rect 8386 9868 8392 9920
rect 8444 9868 8450 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 11348 9908 11376 9948
rect 8996 9880 11376 9908
rect 11532 9908 11560 9948
rect 11882 9936 11888 9988
rect 11940 9936 11946 9988
rect 12434 9936 12440 9988
rect 12492 9936 12498 9988
rect 20892 9979 20950 9985
rect 20892 9945 20904 9979
rect 20938 9976 20950 9979
rect 21266 9976 21272 9988
rect 20938 9948 21272 9976
rect 20938 9945 20950 9948
rect 20892 9939 20950 9945
rect 21266 9936 21272 9948
rect 21324 9936 21330 9988
rect 21358 9936 21364 9988
rect 21416 9976 21422 9988
rect 21910 9976 21916 9988
rect 21416 9948 21916 9976
rect 21416 9936 21422 9948
rect 21910 9936 21916 9948
rect 21968 9976 21974 9988
rect 22281 9979 22339 9985
rect 22281 9976 22293 9979
rect 21968 9948 22293 9976
rect 21968 9936 21974 9948
rect 22281 9945 22293 9948
rect 22327 9945 22339 9979
rect 22664 9976 22692 10007
rect 24412 9976 24440 10007
rect 24578 10004 24584 10056
rect 24636 10004 24642 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 26329 10047 26387 10053
rect 26329 10044 26341 10047
rect 25372 10016 26341 10044
rect 25372 10004 25378 10016
rect 26329 10013 26341 10016
rect 26375 10013 26387 10047
rect 26329 10007 26387 10013
rect 24762 9976 24768 9988
rect 22664 9948 23060 9976
rect 24412 9948 24768 9976
rect 22281 9939 22339 9945
rect 23032 9920 23060 9948
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 24940 9979 24998 9985
rect 24940 9945 24952 9979
rect 24986 9976 24998 9979
rect 24986 9948 26188 9976
rect 24986 9945 24998 9948
rect 24940 9939 24998 9945
rect 12894 9908 12900 9920
rect 11532 9880 12900 9908
rect 8996 9868 9002 9880
rect 12894 9868 12900 9880
rect 12952 9908 12958 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12952 9880 13369 9908
rect 12952 9868 12958 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13357 9871 13415 9877
rect 22094 9868 22100 9920
rect 22152 9868 22158 9920
rect 23014 9868 23020 9920
rect 23072 9908 23078 9920
rect 23109 9911 23167 9917
rect 23109 9908 23121 9911
rect 23072 9880 23121 9908
rect 23072 9868 23078 9880
rect 23109 9877 23121 9880
rect 23155 9877 23167 9911
rect 23109 9871 23167 9877
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9908 24639 9911
rect 25130 9908 25136 9920
rect 24627 9880 25136 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 26050 9868 26056 9920
rect 26108 9868 26114 9920
rect 26160 9917 26188 9948
rect 26145 9911 26203 9917
rect 26145 9877 26157 9911
rect 26191 9877 26203 9911
rect 26145 9871 26203 9877
rect 1104 9818 26864 9840
rect 1104 9766 4829 9818
rect 4881 9766 4893 9818
rect 4945 9766 4957 9818
rect 5009 9766 5021 9818
rect 5073 9766 5085 9818
rect 5137 9766 11268 9818
rect 11320 9766 11332 9818
rect 11384 9766 11396 9818
rect 11448 9766 11460 9818
rect 11512 9766 11524 9818
rect 11576 9766 17707 9818
rect 17759 9766 17771 9818
rect 17823 9766 17835 9818
rect 17887 9766 17899 9818
rect 17951 9766 17963 9818
rect 18015 9766 24146 9818
rect 24198 9766 24210 9818
rect 24262 9766 24274 9818
rect 24326 9766 24338 9818
rect 24390 9766 24402 9818
rect 24454 9766 26864 9818
rect 1104 9744 26864 9766
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4304 9676 4997 9704
rect 4304 9664 4310 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 4985 9667 5043 9673
rect 5810 9664 5816 9716
rect 5868 9664 5874 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6420 9676 7972 9704
rect 6420 9664 6426 9676
rect 7944 9648 7972 9676
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8076 9676 9720 9704
rect 8076 9664 8082 9676
rect 3694 9596 3700 9648
rect 3752 9596 3758 9648
rect 4522 9636 4528 9648
rect 4448 9608 4528 9636
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 4448 9577 4476 9608
rect 4522 9596 4528 9608
rect 4580 9636 4586 9648
rect 5965 9639 6023 9645
rect 5965 9636 5977 9639
rect 4580 9608 5977 9636
rect 4580 9596 4586 9608
rect 5965 9605 5977 9608
rect 6011 9636 6023 9639
rect 6011 9605 6040 9636
rect 5965 9599 6040 9605
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1912 9540 2329 9568
rect 1912 9528 1918 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5224 9540 5549 9568
rect 5224 9528 5230 9540
rect 5537 9537 5549 9540
rect 5583 9568 5595 9571
rect 5810 9568 5816 9580
rect 5583 9540 5816 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6012 9568 6040 9599
rect 6178 9596 6184 9648
rect 6236 9596 6242 9648
rect 6733 9639 6791 9645
rect 6503 9605 6561 9611
rect 6503 9580 6515 9605
rect 6012 9540 6132 9568
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9500 2743 9503
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 2731 9472 4261 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4525 9503 4583 9509
rect 4525 9500 4537 9503
rect 4396 9472 4537 9500
rect 4396 9460 4402 9472
rect 4525 9469 4537 9472
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 5184 9500 5212 9528
rect 4663 9472 5212 9500
rect 5261 9503 5319 9509
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5994 9500 6000 9512
rect 5307 9472 6000 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 4540 9432 4568 9463
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 4540 9404 5304 9432
rect 5276 9376 5304 9404
rect 6104 9376 6132 9540
rect 6454 9528 6460 9580
rect 6512 9571 6515 9580
rect 6549 9602 6561 9605
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 6914 9636 6920 9648
rect 6779 9608 6920 9636
rect 6779 9605 6791 9608
rect 6549 9571 6576 9602
rect 6733 9599 6791 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7834 9596 7840 9648
rect 7892 9596 7898 9648
rect 7926 9596 7932 9648
rect 7984 9596 7990 9648
rect 9306 9636 9312 9648
rect 8496 9608 9312 9636
rect 6512 9568 6576 9571
rect 6512 9540 6583 9568
rect 6512 9528 6518 9540
rect 6555 9500 6583 9540
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7466 9568 7472 9580
rect 7064 9540 7472 9568
rect 7064 9528 7070 9540
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 7742 9568 7748 9580
rect 7699 9540 7748 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8386 9568 8392 9580
rect 8067 9540 8392 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8496 9577 8524 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 8570 9528 8576 9580
rect 8628 9528 8634 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 8938 9568 8944 9580
rect 8803 9540 8944 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9692 9568 9720 9676
rect 21266 9664 21272 9716
rect 21324 9664 21330 9716
rect 21910 9664 21916 9716
rect 21968 9664 21974 9716
rect 22094 9704 22100 9716
rect 22066 9664 22100 9704
rect 22152 9664 22158 9716
rect 24026 9664 24032 9716
rect 24084 9664 24090 9716
rect 25314 9664 25320 9716
rect 25372 9664 25378 9716
rect 10229 9639 10287 9645
rect 10229 9605 10241 9639
rect 10275 9636 10287 9639
rect 10410 9636 10416 9648
rect 10275 9608 10416 9636
rect 10275 9605 10287 9608
rect 10229 9599 10287 9605
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 11609 9639 11667 9645
rect 11609 9605 11621 9639
rect 11655 9636 11667 9639
rect 12434 9636 12440 9648
rect 11655 9608 12440 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 22066 9636 22094 9664
rect 16724 9608 17158 9636
rect 21468 9608 22094 9636
rect 22373 9639 22431 9645
rect 16724 9596 16730 9608
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 9692 9540 10333 9568
rect 10321 9537 10333 9540
rect 10367 9568 10379 9571
rect 11146 9568 11152 9580
rect 10367 9540 11152 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 11146 9528 11152 9540
rect 11204 9568 11210 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 14700 9540 15148 9568
rect 14700 9528 14706 9540
rect 7098 9500 7104 9512
rect 6555 9472 7104 9500
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7374 9460 7380 9512
rect 7432 9460 7438 9512
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 7616 9472 8309 9500
rect 7616 9460 7622 9472
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 8297 9463 8355 9469
rect 15010 9460 15016 9512
rect 15068 9460 15074 9512
rect 15120 9500 15148 9540
rect 18064 9540 18521 9568
rect 18064 9500 18092 9540
rect 18509 9537 18521 9540
rect 18555 9568 18567 9571
rect 19426 9568 19432 9580
rect 18555 9540 19432 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 19426 9528 19432 9540
rect 19484 9528 19490 9580
rect 21468 9577 21496 9608
rect 22373 9605 22385 9639
rect 22419 9636 22431 9639
rect 22922 9636 22928 9648
rect 22419 9608 22928 9636
rect 22419 9605 22431 9608
rect 22373 9599 22431 9605
rect 22922 9596 22928 9608
rect 22980 9636 22986 9648
rect 22980 9608 23152 9636
rect 22980 9596 22986 9608
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 21784 9540 22109 9568
rect 21784 9528 21790 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9568 22615 9571
rect 23014 9568 23020 9580
rect 22603 9540 23020 9568
rect 22603 9537 22615 9540
rect 22557 9531 22615 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 15120 9472 18092 9500
rect 18138 9460 18144 9512
rect 18196 9460 18202 9512
rect 22738 9460 22744 9512
rect 22796 9460 22802 9512
rect 22833 9503 22891 9509
rect 22833 9469 22845 9503
rect 22879 9469 22891 9503
rect 22833 9463 22891 9469
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23124 9500 23152 9608
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 23256 9608 23673 9636
rect 23256 9596 23262 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 23661 9599 23719 9605
rect 23877 9639 23935 9645
rect 23877 9605 23889 9639
rect 23923 9636 23935 9639
rect 24949 9639 25007 9645
rect 23923 9608 24808 9636
rect 23923 9605 23935 9608
rect 23877 9599 23935 9605
rect 24780 9580 24808 9608
rect 24949 9605 24961 9639
rect 24995 9636 25007 9639
rect 25038 9636 25044 9648
rect 24995 9608 25044 9636
rect 24995 9605 25007 9608
rect 24949 9599 25007 9605
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 25165 9639 25223 9645
rect 25165 9605 25177 9639
rect 25211 9636 25223 9639
rect 25777 9639 25835 9645
rect 25777 9636 25789 9639
rect 25211 9608 25789 9636
rect 25211 9605 25223 9608
rect 25165 9599 25223 9605
rect 25777 9605 25789 9608
rect 25823 9605 25835 9639
rect 25777 9599 25835 9605
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 24820 9540 25421 9568
rect 24820 9528 24826 9540
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 26050 9568 26056 9580
rect 25639 9540 26056 9568
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 23382 9500 23388 9512
rect 22971 9472 23388 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 22848 9432 22876 9463
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24578 9460 24584 9512
rect 24636 9500 24642 9512
rect 25608 9500 25636 9531
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 24636 9472 25636 9500
rect 24636 9460 24642 9472
rect 23477 9435 23535 9441
rect 22848 9404 23428 9432
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4111 9367 4169 9373
rect 4111 9364 4123 9367
rect 4028 9336 4123 9364
rect 4028 9324 4034 9336
rect 4111 9333 4123 9336
rect 4157 9364 4169 9367
rect 5166 9364 5172 9376
rect 4157 9336 5172 9364
rect 4157 9333 4169 9336
rect 4111 9327 4169 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5258 9324 5264 9376
rect 5316 9324 5322 9376
rect 5442 9324 5448 9376
rect 5500 9324 5506 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5960 9336 6009 9364
rect 5960 9324 5966 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 5997 9327 6055 9333
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6144 9336 6377 9364
rect 6144 9324 6150 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 7006 9364 7012 9376
rect 6595 9336 7012 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9364 8263 9367
rect 11882 9364 11888 9376
rect 8251 9336 11888 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 13814 9364 13820 9376
rect 12860 9336 13820 9364
rect 12860 9324 12866 9336
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 16439 9367 16497 9373
rect 16439 9364 16451 9367
rect 15804 9336 16451 9364
rect 15804 9324 15810 9336
rect 16439 9333 16451 9336
rect 16485 9333 16497 9367
rect 16439 9327 16497 9333
rect 16758 9324 16764 9376
rect 16816 9324 16822 9376
rect 22186 9324 22192 9376
rect 22244 9324 22250 9376
rect 23198 9324 23204 9376
rect 23256 9324 23262 9376
rect 23400 9364 23428 9404
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 23934 9432 23940 9444
rect 23523 9404 23940 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 23934 9392 23940 9404
rect 23992 9392 23998 9444
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23400 9336 23857 9364
rect 23845 9333 23857 9336
rect 23891 9364 23903 9367
rect 24578 9364 24584 9376
rect 23891 9336 24584 9364
rect 23891 9333 23903 9336
rect 23845 9327 23903 9333
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 25130 9324 25136 9376
rect 25188 9324 25194 9376
rect 1104 9274 26864 9296
rect 1104 9222 4169 9274
rect 4221 9222 4233 9274
rect 4285 9222 4297 9274
rect 4349 9222 4361 9274
rect 4413 9222 4425 9274
rect 4477 9222 10608 9274
rect 10660 9222 10672 9274
rect 10724 9222 10736 9274
rect 10788 9222 10800 9274
rect 10852 9222 10864 9274
rect 10916 9222 17047 9274
rect 17099 9222 17111 9274
rect 17163 9222 17175 9274
rect 17227 9222 17239 9274
rect 17291 9222 17303 9274
rect 17355 9222 23486 9274
rect 23538 9222 23550 9274
rect 23602 9222 23614 9274
rect 23666 9222 23678 9274
rect 23730 9222 23742 9274
rect 23794 9222 26864 9274
rect 1104 9200 26864 9222
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 2866 9160 2872 9172
rect 2823 9132 2872 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 5994 9120 6000 9172
rect 6052 9120 6058 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7156 9132 7481 9160
rect 7156 9120 7162 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 10965 9163 11023 9169
rect 10965 9129 10977 9163
rect 11011 9160 11023 9163
rect 11054 9160 11060 9172
rect 11011 9132 11060 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12575 9132 13001 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 4341 9095 4399 9101
rect 4341 9061 4353 9095
rect 4387 9092 4399 9095
rect 4614 9092 4620 9104
rect 4387 9064 4620 9092
rect 4387 9061 4399 9064
rect 4341 9055 4399 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 6178 9092 6184 9104
rect 5500 9064 6184 9092
rect 5500 9052 5506 9064
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 12345 9095 12403 9101
rect 6288 9064 8800 9092
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6288 9024 6316 9064
rect 5960 8996 6316 9024
rect 7837 9027 7895 9033
rect 5960 8984 5966 8996
rect 7837 8993 7849 9027
rect 7883 9024 7895 9027
rect 8662 9024 8668 9036
rect 7883 8996 8668 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 8772 9024 8800 9064
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 12802 9092 12808 9104
rect 12391 9064 12808 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 13004 9092 13032 9123
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 13136 9132 13461 9160
rect 13136 9120 13142 9132
rect 13449 9129 13461 9132
rect 13495 9160 13507 9163
rect 13722 9160 13728 9172
rect 13495 9132 13728 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 13722 9120 13728 9132
rect 13780 9160 13786 9172
rect 14090 9160 14096 9172
rect 13780 9132 14096 9160
rect 13780 9120 13786 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15620 9132 15669 9160
rect 15620 9120 15626 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 17497 9163 17555 9169
rect 17497 9129 17509 9163
rect 17543 9160 17555 9163
rect 18138 9160 18144 9172
rect 17543 9132 18144 9160
rect 17543 9129 17555 9132
rect 17497 9123 17555 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18472 9132 18889 9160
rect 18472 9120 18478 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 21729 9163 21787 9169
rect 21729 9129 21741 9163
rect 21775 9160 21787 9163
rect 22186 9160 22192 9172
rect 21775 9132 22192 9160
rect 21775 9129 21787 9132
rect 21729 9123 21787 9129
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23256 9132 23673 9160
rect 23256 9120 23262 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 13630 9092 13636 9104
rect 13004 9064 13636 9092
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 17405 9095 17463 9101
rect 17405 9061 17417 9095
rect 17451 9092 17463 9095
rect 19242 9092 19248 9104
rect 17451 9064 18184 9092
rect 17451 9061 17463 9064
rect 17405 9055 17463 9061
rect 8772 8996 13400 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 2958 8956 2964 8968
rect 2915 8928 2964 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 5920 8956 5948 8984
rect 4019 8928 5948 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 12728 8928 13216 8956
rect 7668 8888 7696 8919
rect 7668 8860 8616 8888
rect 8588 8832 8616 8860
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10778 8888 10784 8900
rect 10192 8860 10784 8888
rect 10192 8848 10198 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 12728 8897 12756 8928
rect 13188 8900 13216 8928
rect 12497 8891 12555 8897
rect 12497 8888 12509 8891
rect 11756 8860 12509 8888
rect 11756 8848 11762 8860
rect 12497 8857 12509 8860
rect 12543 8857 12555 8891
rect 12497 8851 12555 8857
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8857 12771 8891
rect 12713 8851 12771 8857
rect 12894 8848 12900 8900
rect 12952 8897 12958 8900
rect 12952 8891 13015 8897
rect 12952 8857 12969 8891
rect 13003 8857 13015 8891
rect 12952 8851 13015 8857
rect 12952 8848 12958 8851
rect 13170 8848 13176 8900
rect 13228 8848 13234 8900
rect 13262 8848 13268 8900
rect 13320 8848 13326 8900
rect 13372 8888 13400 8996
rect 17126 8984 17132 9036
rect 17184 8984 17190 9036
rect 18046 9024 18052 9036
rect 17696 8996 18052 9024
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 16022 8956 16028 8968
rect 15611 8928 16028 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 13465 8891 13523 8897
rect 13465 8888 13477 8891
rect 13372 8860 13477 8888
rect 13465 8857 13477 8860
rect 13511 8857 13523 8891
rect 13465 8851 13523 8857
rect 15378 8848 15384 8900
rect 15436 8888 15442 8900
rect 16592 8888 16620 8919
rect 16758 8916 16764 8968
rect 16816 8956 16822 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16816 8928 17049 8956
rect 16816 8916 16822 8928
rect 17037 8925 17049 8928
rect 17083 8956 17095 8959
rect 17218 8956 17224 8968
rect 17083 8928 17224 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17696 8965 17724 8996
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 18156 9033 18184 9064
rect 18892 9064 19248 9092
rect 18141 9027 18199 9033
rect 18141 8993 18153 9027
rect 18187 8993 18199 9027
rect 18141 8987 18199 8993
rect 18230 8984 18236 9036
rect 18288 8984 18294 9036
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8956 17923 8959
rect 18892 8956 18920 9064
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 19426 9052 19432 9104
rect 19484 9092 19490 9104
rect 19484 9064 22048 9092
rect 19484 9052 19490 9064
rect 21818 9024 21824 9036
rect 20640 8996 21824 9024
rect 20640 8965 20668 8996
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22020 9033 22048 9064
rect 23290 9052 23296 9104
rect 23348 9092 23354 9104
rect 23477 9095 23535 9101
rect 23477 9092 23489 9095
rect 23348 9064 23489 9092
rect 23348 9052 23354 9064
rect 23477 9061 23489 9064
rect 23523 9061 23535 9095
rect 23477 9055 23535 9061
rect 24026 9052 24032 9104
rect 24084 9052 24090 9104
rect 22005 9027 22063 9033
rect 22005 8993 22017 9027
rect 22051 8993 22063 9027
rect 24486 9024 24492 9036
rect 22005 8987 22063 8993
rect 23952 8996 24492 9024
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 17911 8928 18920 8956
rect 18984 8928 19441 8956
rect 17911 8925 17923 8928
rect 17865 8919 17923 8925
rect 15436 8860 16620 8888
rect 17773 8891 17831 8897
rect 15436 8848 15442 8860
rect 17773 8857 17785 8891
rect 17819 8857 17831 8891
rect 17773 8851 17831 8857
rect 18003 8891 18061 8897
rect 18003 8857 18015 8891
rect 18049 8888 18061 8891
rect 18049 8860 18276 8888
rect 18049 8857 18061 8860
rect 18003 8851 18061 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2130 8820 2136 8832
rect 1627 8792 2136 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 10981 8823 11039 8829
rect 10981 8820 10993 8823
rect 8628 8792 10993 8820
rect 8628 8780 8634 8792
rect 10981 8789 10993 8792
rect 11027 8789 11039 8823
rect 10981 8783 11039 8789
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 12066 8820 12072 8832
rect 11195 8792 12072 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12802 8780 12808 8832
rect 12860 8780 12866 8832
rect 13633 8823 13691 8829
rect 13633 8789 13645 8823
rect 13679 8820 13691 8823
rect 15102 8820 15108 8832
rect 13679 8792 15108 8820
rect 13679 8789 13691 8792
rect 13633 8783 13691 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 17788 8820 17816 8851
rect 18138 8820 18144 8832
rect 17788 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18248 8820 18276 8860
rect 18414 8848 18420 8900
rect 18472 8848 18478 8900
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8857 18659 8891
rect 18601 8851 18659 8857
rect 18322 8820 18328 8832
rect 18248 8792 18328 8820
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 18616 8820 18644 8851
rect 18690 8848 18696 8900
rect 18748 8848 18754 8900
rect 18898 8891 18956 8897
rect 18898 8888 18910 8891
rect 18800 8860 18910 8888
rect 18800 8820 18828 8860
rect 18898 8857 18910 8860
rect 18944 8888 18956 8891
rect 18984 8888 19012 8928
rect 19429 8925 19441 8928
rect 19475 8956 19487 8959
rect 20625 8959 20683 8965
rect 19475 8928 20484 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 20346 8888 20352 8900
rect 18944 8860 19012 8888
rect 19076 8860 20352 8888
rect 18944 8857 18956 8860
rect 18898 8851 18956 8857
rect 19076 8829 19104 8860
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 20456 8888 20484 8928
rect 20625 8925 20637 8959
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8925 21419 8959
rect 22020 8956 22048 8987
rect 23952 8956 23980 8996
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 22020 8928 23980 8956
rect 25777 8959 25835 8965
rect 21361 8919 21419 8925
rect 25777 8925 25789 8959
rect 25823 8956 25835 8959
rect 26326 8956 26332 8968
rect 25823 8928 26332 8956
rect 25823 8925 25835 8928
rect 25777 8919 25835 8925
rect 21266 8888 21272 8900
rect 20456 8860 21272 8888
rect 21266 8848 21272 8860
rect 21324 8848 21330 8900
rect 21376 8888 21404 8919
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 22094 8888 22100 8900
rect 21376 8860 22100 8888
rect 22094 8848 22100 8860
rect 22152 8848 22158 8900
rect 22272 8891 22330 8897
rect 22272 8857 22284 8891
rect 22318 8888 22330 8891
rect 22462 8888 22468 8900
rect 22318 8860 22468 8888
rect 22318 8857 22330 8860
rect 22272 8851 22330 8857
rect 22462 8848 22468 8860
rect 22520 8848 22526 8900
rect 18564 8792 18828 8820
rect 19061 8823 19119 8829
rect 18564 8780 18570 8792
rect 19061 8789 19073 8823
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 19334 8780 19340 8832
rect 19392 8780 19398 8832
rect 20530 8780 20536 8832
rect 20588 8780 20594 8832
rect 21726 8780 21732 8832
rect 21784 8780 21790 8832
rect 21913 8823 21971 8829
rect 21913 8789 21925 8823
rect 21959 8820 21971 8823
rect 22646 8820 22652 8832
rect 21959 8792 22652 8820
rect 21959 8789 21971 8792
rect 21913 8783 21971 8789
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 23382 8780 23388 8832
rect 23440 8780 23446 8832
rect 23658 8780 23664 8832
rect 23716 8780 23722 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 1104 8730 26864 8752
rect 1104 8678 4829 8730
rect 4881 8678 4893 8730
rect 4945 8678 4957 8730
rect 5009 8678 5021 8730
rect 5073 8678 5085 8730
rect 5137 8678 11268 8730
rect 11320 8678 11332 8730
rect 11384 8678 11396 8730
rect 11448 8678 11460 8730
rect 11512 8678 11524 8730
rect 11576 8678 17707 8730
rect 17759 8678 17771 8730
rect 17823 8678 17835 8730
rect 17887 8678 17899 8730
rect 17951 8678 17963 8730
rect 18015 8678 24146 8730
rect 24198 8678 24210 8730
rect 24262 8678 24274 8730
rect 24326 8678 24338 8730
rect 24390 8678 24402 8730
rect 24454 8678 26864 8730
rect 1104 8656 26864 8678
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 8731 8619 8789 8625
rect 8731 8616 8743 8619
rect 6236 8588 8743 8616
rect 6236 8576 6242 8588
rect 8731 8585 8743 8588
rect 8777 8585 8789 8619
rect 8731 8579 8789 8585
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13228 8588 13645 8616
rect 13228 8576 13234 8588
rect 13633 8585 13645 8588
rect 13679 8616 13691 8619
rect 13722 8616 13728 8628
rect 13679 8588 13728 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 13722 8576 13728 8588
rect 13780 8616 13786 8628
rect 14182 8616 14188 8628
rect 13780 8588 14188 8616
rect 13780 8576 13786 8588
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 15068 8588 17141 8616
rect 15068 8576 15074 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17368 8588 18184 8616
rect 17368 8576 17374 8588
rect 8941 8551 8999 8557
rect 8941 8517 8953 8551
rect 8987 8548 8999 8551
rect 9122 8548 9128 8560
rect 8987 8520 9128 8548
rect 8987 8517 8999 8520
rect 8941 8511 8999 8517
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 13357 8551 13415 8557
rect 13357 8548 13369 8551
rect 12860 8520 13369 8548
rect 12860 8508 12866 8520
rect 13357 8517 13369 8520
rect 13403 8517 13415 8551
rect 13357 8511 13415 8517
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 13504 8520 14105 8548
rect 13504 8508 13510 8520
rect 14093 8517 14105 8520
rect 14139 8548 14151 8551
rect 14458 8548 14464 8560
rect 14139 8520 14464 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 15746 8508 15752 8560
rect 15804 8548 15810 8560
rect 18156 8548 18184 8588
rect 18322 8576 18328 8628
rect 18380 8616 18386 8628
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 18380 8588 18429 8616
rect 18380 8576 18386 8588
rect 18417 8585 18429 8588
rect 18463 8616 18475 8619
rect 19518 8616 19524 8628
rect 18463 8588 19524 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 22462 8576 22468 8628
rect 22520 8576 22526 8628
rect 22738 8576 22744 8628
rect 22796 8576 22802 8628
rect 23934 8616 23940 8628
rect 23860 8588 23940 8616
rect 18506 8548 18512 8560
rect 15804 8520 18092 8548
rect 18156 8520 18512 8548
rect 15804 8508 15810 8520
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 9030 8480 9036 8492
rect 5592 8452 9036 8480
rect 5592 8440 5598 8452
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 13078 8440 13084 8492
rect 13136 8480 13142 8492
rect 13136 8452 13584 8480
rect 13136 8440 13142 8452
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 8444 8316 8585 8344
rect 8444 8304 8450 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 8573 8307 8631 8313
rect 12894 8304 12900 8356
rect 12952 8304 12958 8356
rect 13280 8344 13308 8375
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 13280 8316 13461 8344
rect 13449 8313 13461 8316
rect 13495 8313 13507 8347
rect 13556 8344 13584 8452
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13688 8452 14013 8480
rect 13688 8440 13694 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15286 8480 15292 8492
rect 15243 8452 15292 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17184 8452 17908 8480
rect 17184 8440 17190 8452
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14148 8384 14412 8412
rect 14148 8372 14154 8384
rect 14384 8353 14412 8384
rect 15378 8372 15384 8424
rect 15436 8372 15442 8424
rect 17310 8372 17316 8424
rect 17368 8372 17374 8424
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17589 8415 17647 8421
rect 17589 8381 17601 8415
rect 17635 8412 17647 8415
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 17635 8384 17785 8412
rect 17635 8381 17647 8384
rect 17589 8375 17647 8381
rect 17773 8381 17785 8384
rect 17819 8381 17831 8415
rect 17880 8412 17908 8452
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 18064 8480 18092 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 20530 8508 20536 8560
rect 20588 8508 20594 8560
rect 23658 8548 23664 8560
rect 22066 8520 23664 8548
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18064 8452 18245 8480
rect 18233 8449 18245 8452
rect 18279 8480 18291 8483
rect 18322 8480 18328 8492
rect 18279 8452 18328 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18322 8440 18328 8452
rect 18380 8480 18386 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 18380 8452 18613 8480
rect 18380 8440 18386 8452
rect 18601 8449 18613 8452
rect 18647 8480 18659 8483
rect 18690 8480 18696 8492
rect 18647 8452 18696 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18923 8452 19165 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 19153 8443 19211 8449
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17880 8384 18153 8412
rect 17773 8375 17831 8381
rect 18141 8381 18153 8384
rect 18187 8412 18199 8415
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18187 8384 18797 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 18785 8381 18797 8384
rect 18831 8412 18843 8415
rect 18966 8412 18972 8424
rect 18831 8384 18972 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 14369 8347 14427 8353
rect 13556 8316 14044 8344
rect 13449 8307 13507 8313
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 9766 8276 9772 8288
rect 8803 8248 9772 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 13354 8236 13360 8288
rect 13412 8236 13418 8288
rect 13633 8279 13691 8285
rect 13633 8245 13645 8279
rect 13679 8276 13691 8279
rect 13906 8276 13912 8288
rect 13679 8248 13912 8276
rect 13679 8245 13691 8248
rect 13633 8239 13691 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14016 8276 14044 8316
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 17218 8344 17224 8356
rect 15068 8316 17224 8344
rect 15068 8304 15074 8316
rect 17218 8304 17224 8316
rect 17276 8344 17282 8356
rect 17512 8344 17540 8375
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19260 8412 19288 8443
rect 19426 8440 19432 8492
rect 19484 8440 19490 8492
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 21726 8480 21732 8492
rect 20772 8452 21732 8480
rect 20772 8440 20778 8452
rect 21726 8440 21732 8452
rect 21784 8480 21790 8492
rect 22066 8480 22094 8520
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 23860 8557 23888 8588
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 23854 8551 23912 8557
rect 23854 8517 23866 8551
rect 23900 8517 23912 8551
rect 23854 8511 23912 8517
rect 21784 8452 22094 8480
rect 21784 8440 21790 8452
rect 22646 8440 22652 8492
rect 22704 8440 22710 8492
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8480 24179 8483
rect 24486 8480 24492 8492
rect 24167 8452 24492 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 24486 8440 24492 8452
rect 24544 8440 24550 8492
rect 19116 8384 19288 8412
rect 19116 8372 19122 8384
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 17954 8344 17960 8356
rect 17276 8316 17960 8344
rect 17276 8304 17282 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18046 8304 18052 8356
rect 18104 8304 18110 8356
rect 18690 8344 18696 8356
rect 18432 8316 18696 8344
rect 14090 8276 14096 8288
rect 14016 8248 14096 8276
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 14553 8279 14611 8285
rect 14553 8245 14565 8279
rect 14599 8276 14611 8279
rect 14826 8276 14832 8288
rect 14599 8248 14832 8276
rect 14599 8245 14611 8248
rect 14553 8239 14611 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 17972 8276 18000 8304
rect 18432 8288 18460 8316
rect 18690 8304 18696 8316
rect 18748 8304 18754 8356
rect 18414 8276 18420 8288
rect 17972 8248 18420 8276
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 21223 8279 21281 8285
rect 21223 8276 21235 8279
rect 20036 8248 21235 8276
rect 20036 8236 20042 8248
rect 21223 8245 21235 8248
rect 21269 8276 21281 8279
rect 21634 8276 21640 8288
rect 21269 8248 21640 8276
rect 21269 8245 21281 8248
rect 21223 8239 21281 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 1104 8186 26864 8208
rect 1104 8134 4169 8186
rect 4221 8134 4233 8186
rect 4285 8134 4297 8186
rect 4349 8134 4361 8186
rect 4413 8134 4425 8186
rect 4477 8134 10608 8186
rect 10660 8134 10672 8186
rect 10724 8134 10736 8186
rect 10788 8134 10800 8186
rect 10852 8134 10864 8186
rect 10916 8134 17047 8186
rect 17099 8134 17111 8186
rect 17163 8134 17175 8186
rect 17227 8134 17239 8186
rect 17291 8134 17303 8186
rect 17355 8134 23486 8186
rect 23538 8134 23550 8186
rect 23602 8134 23614 8186
rect 23666 8134 23678 8186
rect 23730 8134 23742 8186
rect 23794 8134 26864 8186
rect 1104 8112 26864 8134
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 12032 8044 12081 8072
rect 12032 8032 12038 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 12986 8072 12992 8084
rect 12851 8044 12992 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13630 8072 13636 8084
rect 13587 8044 13636 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14148 8044 15884 8072
rect 14148 8032 14154 8044
rect 10962 7964 10968 8016
rect 11020 8004 11026 8016
rect 11057 8007 11115 8013
rect 11057 8004 11069 8007
rect 11020 7976 11069 8004
rect 11020 7964 11026 7976
rect 11057 7973 11069 7976
rect 11103 7973 11115 8007
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 11057 7967 11115 7973
rect 12268 7976 12633 8004
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 4065 7939 4123 7945
rect 2271 7908 2774 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2130 7828 2136 7880
rect 2188 7828 2194 7880
rect 2746 7800 2774 7908
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 5626 7936 5632 7948
rect 4111 7908 5632 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 9582 7936 9588 7948
rect 7024 7908 9588 7936
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4246 7828 4252 7880
rect 4304 7828 4310 7880
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4522 7868 4528 7880
rect 4387 7840 4528 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 7024 7877 7052 7908
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 12268 7945 12296 7976
rect 12621 7973 12633 7976
rect 12667 7973 12679 8007
rect 12621 7967 12679 7973
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 12768 7976 14473 8004
rect 12768 7964 12774 7976
rect 14461 7973 14473 7976
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 12253 7939 12311 7945
rect 11348 7908 11652 7936
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7248 7840 7573 7868
rect 7248 7828 7254 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8294 7868 8300 7880
rect 7975 7840 8300 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10134 7868 10140 7880
rect 9180 7840 10140 7868
rect 9180 7828 9186 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 11348 7877 11376 7908
rect 11624 7877 11652 7908
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13446 7936 13452 7948
rect 13219 7908 13452 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 13909 7939 13967 7945
rect 13909 7936 13921 7939
rect 13780 7908 13921 7936
rect 13780 7896 13786 7908
rect 13909 7905 13921 7908
rect 13955 7936 13967 7939
rect 13955 7908 14320 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11882 7868 11888 7880
rect 11655 7840 11888 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 2746 7772 7420 7800
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3844 7704 3893 7732
rect 3844 7692 3850 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 7392 7732 7420 7772
rect 7466 7760 7472 7812
rect 7524 7800 7530 7812
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 7524 7772 7757 7800
rect 7524 7760 7530 7772
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 7745 7763 7803 7769
rect 7837 7803 7895 7809
rect 7837 7769 7849 7803
rect 7883 7769 7895 7803
rect 7837 7763 7895 7769
rect 7852 7732 7880 7763
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 8260 7772 8953 7800
rect 8260 7760 8266 7772
rect 8941 7769 8953 7772
rect 8987 7769 8999 7803
rect 8941 7763 8999 7769
rect 9309 7803 9367 7809
rect 9309 7769 9321 7803
rect 9355 7800 9367 7803
rect 9766 7800 9772 7812
rect 9355 7772 9772 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 9766 7760 9772 7772
rect 9824 7800 9830 7812
rect 10686 7800 10692 7812
rect 9824 7772 10692 7800
rect 9824 7760 9830 7772
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 11054 7760 11060 7812
rect 11112 7760 11118 7812
rect 11241 7803 11299 7809
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 11440 7800 11468 7831
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 13078 7868 13084 7880
rect 12391 7840 13084 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 14292 7877 14320 7908
rect 14844 7908 15240 7936
rect 14642 7877 14648 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13688 7840 14105 7868
rect 13688 7828 13694 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14640 7831 14648 7877
rect 14700 7868 14706 7880
rect 14844 7868 14872 7908
rect 14700 7840 14872 7868
rect 14642 7828 14648 7831
rect 14700 7828 14706 7840
rect 15010 7828 15016 7880
rect 15068 7828 15074 7880
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 15212 7868 15240 7908
rect 15335 7871 15393 7877
rect 15335 7868 15347 7871
rect 15212 7840 15347 7868
rect 15335 7837 15347 7840
rect 15381 7837 15393 7871
rect 15335 7831 15393 7837
rect 15746 7828 15752 7880
rect 15804 7828 15810 7880
rect 15856 7877 15884 8044
rect 18138 8032 18144 8084
rect 18196 8032 18202 8084
rect 18322 8032 18328 8084
rect 18380 8032 18386 8084
rect 19794 8032 19800 8084
rect 19852 8032 19858 8084
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20404 8044 20944 8072
rect 20404 8032 20410 8044
rect 19334 8004 19340 8016
rect 18432 7976 19340 8004
rect 18432 7945 18460 7976
rect 19334 7964 19340 7976
rect 19392 8004 19398 8016
rect 20806 8004 20812 8016
rect 19392 7976 20812 8004
rect 19392 7964 19398 7976
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7905 18475 7939
rect 18417 7899 18475 7905
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 18923 7908 19656 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 18966 7828 18972 7880
rect 19024 7828 19030 7880
rect 19242 7828 19248 7880
rect 19300 7828 19306 7880
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19628 7877 19656 7908
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 19944 7908 19993 7936
rect 19944 7896 19950 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 20070 7896 20076 7948
rect 20128 7896 20134 7948
rect 20165 7939 20223 7945
rect 20165 7905 20177 7939
rect 20211 7936 20223 7939
rect 20438 7936 20444 7948
rect 20211 7908 20444 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 20622 7936 20628 7948
rect 20548 7908 20628 7936
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 20254 7828 20260 7880
rect 20312 7828 20318 7880
rect 20548 7877 20576 7908
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20916 7868 20944 8044
rect 20990 7868 20996 7880
rect 20763 7840 20996 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 11698 7800 11704 7812
rect 11287 7772 11704 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 13541 7803 13599 7809
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14458 7800 14464 7812
rect 13587 7772 14464 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 14734 7760 14740 7812
rect 14792 7760 14798 7812
rect 14826 7760 14832 7812
rect 14884 7800 14890 7812
rect 14884 7772 15424 7800
rect 14884 7760 14890 7772
rect 8018 7732 8024 7744
rect 7392 7704 8024 7732
rect 3881 7695 3939 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8754 7732 8760 7744
rect 8159 7704 8760 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 11517 7735 11575 7741
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 11606 7732 11612 7744
rect 11563 7704 11612 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12492 7704 12541 7732
rect 12492 7692 12498 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 15102 7732 15108 7744
rect 12851 7704 15108 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 15194 7692 15200 7744
rect 15252 7692 15258 7744
rect 15396 7732 15424 7772
rect 15470 7760 15476 7812
rect 15528 7760 15534 7812
rect 15565 7803 15623 7809
rect 15565 7769 15577 7803
rect 15611 7769 15623 7803
rect 15565 7763 15623 7769
rect 19429 7803 19487 7809
rect 19429 7769 19441 7803
rect 19475 7800 19487 7803
rect 19794 7800 19800 7812
rect 19475 7772 19800 7800
rect 19475 7769 19487 7772
rect 19429 7763 19487 7769
rect 15580 7732 15608 7763
rect 19794 7760 19800 7772
rect 19852 7760 19858 7812
rect 15396 7704 15608 7732
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 19886 7732 19892 7744
rect 18196 7704 19892 7732
rect 18196 7692 18202 7704
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 20622 7732 20628 7744
rect 20487 7704 20628 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 20898 7692 20904 7744
rect 20956 7692 20962 7744
rect 1104 7642 26864 7664
rect 1104 7590 4829 7642
rect 4881 7590 4893 7642
rect 4945 7590 4957 7642
rect 5009 7590 5021 7642
rect 5073 7590 5085 7642
rect 5137 7590 11268 7642
rect 11320 7590 11332 7642
rect 11384 7590 11396 7642
rect 11448 7590 11460 7642
rect 11512 7590 11524 7642
rect 11576 7590 17707 7642
rect 17759 7590 17771 7642
rect 17823 7590 17835 7642
rect 17887 7590 17899 7642
rect 17951 7590 17963 7642
rect 18015 7590 24146 7642
rect 24198 7590 24210 7642
rect 24262 7590 24274 7642
rect 24326 7590 24338 7642
rect 24390 7590 24402 7642
rect 24454 7590 26864 7642
rect 1104 7568 26864 7590
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4304 7500 4537 7528
rect 4304 7488 4310 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 7466 7488 7472 7540
rect 7524 7488 7530 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 7975 7500 11836 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 3510 7420 3516 7472
rect 3568 7420 3574 7472
rect 5626 7420 5632 7472
rect 5684 7420 5690 7472
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3421 7395 3479 7401
rect 3421 7392 3433 7395
rect 3191 7364 3433 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3421 7361 3433 7364
rect 3467 7361 3479 7395
rect 3528 7392 3556 7420
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3528 7364 3709 7392
rect 3421 7355 3479 7361
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4614 7392 4620 7404
rect 4019 7364 4620 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 3436 7324 3464 7355
rect 3878 7324 3884 7336
rect 3436 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3988 7256 4016 7355
rect 4614 7352 4620 7364
rect 4672 7392 4678 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4672 7364 4997 7392
rect 4672 7352 4678 7364
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5350 7392 5356 7404
rect 5031 7364 5356 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5350 7352 5356 7364
rect 5408 7392 5414 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5408 7364 5457 7392
rect 5408 7352 5414 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5166 7324 5172 7336
rect 5123 7296 5172 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5460 7324 5488 7355
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7484 7392 7512 7488
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8076 7432 8493 7460
rect 8076 7420 8082 7432
rect 8481 7429 8493 7432
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 8754 7420 8760 7472
rect 8812 7420 8818 7472
rect 11808 7460 11836 7500
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 12710 7528 12716 7540
rect 12084 7500 12716 7528
rect 12084 7460 12112 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13357 7531 13415 7537
rect 13357 7497 13369 7531
rect 13403 7528 13415 7531
rect 13722 7528 13728 7540
rect 13403 7500 13728 7528
rect 13403 7497 13415 7500
rect 13357 7491 13415 7497
rect 13722 7488 13728 7500
rect 13780 7528 13786 7540
rect 14182 7528 14188 7540
rect 13780 7500 14188 7528
rect 13780 7488 13786 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14642 7488 14648 7540
rect 14700 7528 14706 7540
rect 14737 7531 14795 7537
rect 14737 7528 14749 7531
rect 14700 7500 14749 7528
rect 14700 7488 14706 7500
rect 14737 7497 14749 7500
rect 14783 7497 14795 7531
rect 14737 7491 14795 7497
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 17000 7500 17233 7528
rect 17000 7488 17006 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 17221 7491 17279 7497
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 18782 7528 18788 7540
rect 17911 7500 18788 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 19484 7500 19533 7528
rect 19484 7488 19490 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 19521 7491 19579 7497
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 19852 7500 21189 7528
rect 19852 7488 19858 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 9048 7432 9720 7460
rect 7423 7364 7512 7392
rect 7837 7395 7895 7401
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 7852 7324 7880 7355
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8711 7364 8861 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8849 7361 8861 7364
rect 8895 7392 8907 7395
rect 8938 7392 8944 7404
rect 8895 7364 8944 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 5460 7296 7880 7324
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 9048 7324 9076 7432
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9692 7401 9720 7432
rect 11256 7432 11652 7460
rect 11808 7432 12112 7460
rect 12161 7463 12219 7469
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 8588 7296 9076 7324
rect 3292 7228 4016 7256
rect 3292 7216 3298 7228
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 8588 7256 8616 7296
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 10042 7324 10048 7336
rect 9539 7296 10048 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10134 7284 10140 7336
rect 10192 7284 10198 7336
rect 10594 7333 10600 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10244 7296 10425 7324
rect 7340 7228 8616 7256
rect 7340 7216 7346 7228
rect 8662 7216 8668 7268
rect 8720 7256 8726 7268
rect 10244 7256 10272 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10551 7327 10600 7333
rect 10551 7293 10563 7327
rect 10597 7293 10600 7327
rect 10551 7287 10600 7293
rect 10594 7284 10600 7287
rect 10652 7284 10658 7336
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11256 7324 11284 7432
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10744 7296 11284 7324
rect 11348 7364 11529 7392
rect 10744 7284 10750 7296
rect 8720 7228 10272 7256
rect 8720 7216 8726 7228
rect 3050 7148 3056 7200
rect 3108 7148 3114 7200
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4856 7160 5273 7188
rect 4856 7148 4862 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 5902 7188 5908 7200
rect 5859 7160 5908 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 9122 7188 9128 7200
rect 7423 7160 9128 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9766 7188 9772 7200
rect 9447 7160 9772 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11348 7197 11376 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11624 7324 11652 7432
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 13446 7460 13452 7472
rect 12207 7432 13452 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 13817 7463 13875 7469
rect 13817 7429 13829 7463
rect 13863 7429 13875 7463
rect 13817 7423 13875 7429
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 11790 7392 11796 7404
rect 11747 7364 11796 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13630 7392 13636 7404
rect 13035 7364 13636 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13832 7392 13860 7423
rect 13998 7420 14004 7472
rect 14056 7460 14062 7472
rect 14277 7463 14335 7469
rect 14277 7460 14289 7463
rect 14056 7432 14289 7460
rect 14056 7420 14062 7432
rect 14277 7429 14289 7432
rect 14323 7429 14335 7463
rect 19978 7460 19984 7472
rect 14277 7423 14335 7429
rect 17696 7432 19984 7460
rect 17696 7404 17724 7432
rect 19978 7420 19984 7432
rect 20036 7420 20042 7472
rect 20257 7463 20315 7469
rect 20257 7429 20269 7463
rect 20303 7460 20315 7463
rect 20898 7460 20904 7472
rect 20303 7432 20904 7460
rect 20303 7429 20315 7432
rect 20257 7423 20315 7429
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 21082 7420 21088 7472
rect 21140 7460 21146 7472
rect 21421 7463 21479 7469
rect 21421 7460 21433 7463
rect 21140 7432 21433 7460
rect 21140 7420 21146 7432
rect 21421 7429 21433 7432
rect 21467 7429 21479 7463
rect 21421 7423 21479 7429
rect 21634 7420 21640 7472
rect 21692 7420 21698 7472
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 13832 7364 16773 7392
rect 16761 7361 16773 7364
rect 16807 7392 16819 7395
rect 16942 7392 16948 7404
rect 16807 7364 16948 7392
rect 16807 7361 16819 7364
rect 16761 7355 16819 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17092 7364 17417 7392
rect 17092 7352 17098 7364
rect 17405 7361 17417 7364
rect 17451 7392 17463 7395
rect 17678 7392 17684 7404
rect 17451 7364 17684 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 18138 7392 18144 7404
rect 17911 7364 18144 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 11624 7296 12572 7324
rect 12544 7265 12572 7296
rect 12529 7259 12587 7265
rect 12529 7225 12541 7259
rect 12575 7256 12587 7259
rect 12986 7256 12992 7268
rect 12575 7228 12992 7256
rect 12575 7225 12587 7228
rect 12529 7219 12587 7225
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 13648 7256 13676 7352
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 16853 7327 16911 7333
rect 14516 7296 16712 7324
rect 14516 7284 14522 7296
rect 13648 7228 13860 7256
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11204 7160 11345 7188
rect 11204 7148 11210 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 12158 7148 12164 7200
rect 12216 7148 12222 7200
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13446 7188 13452 7200
rect 13403 7160 13452 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13538 7148 13544 7200
rect 13596 7148 13602 7200
rect 13630 7148 13636 7200
rect 13688 7148 13694 7200
rect 13832 7197 13860 7228
rect 14182 7216 14188 7268
rect 14240 7216 14246 7268
rect 14550 7216 14556 7268
rect 14608 7216 14614 7268
rect 16684 7256 16712 7296
rect 16853 7293 16865 7327
rect 16899 7324 16911 7327
rect 17880 7324 17908 7355
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 20070 7392 20076 7404
rect 19300 7364 20076 7392
rect 19300 7352 19306 7364
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 16899 7296 17908 7324
rect 16899 7293 16911 7296
rect 16853 7287 16911 7293
rect 16868 7256 16896 7287
rect 19518 7284 19524 7336
rect 19576 7324 19582 7336
rect 20364 7324 20392 7355
rect 19576 7296 20392 7324
rect 20456 7324 20484 7355
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20680 7364 20729 7392
rect 20680 7352 20686 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 20990 7352 20996 7404
rect 21048 7352 21054 7404
rect 20898 7324 20904 7336
rect 20456 7296 20904 7324
rect 19576 7284 19582 7296
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 16684 7228 16896 7256
rect 16942 7216 16948 7268
rect 17000 7256 17006 7268
rect 17681 7259 17739 7265
rect 17681 7256 17693 7259
rect 17000 7228 17693 7256
rect 17000 7216 17006 7228
rect 17681 7225 17693 7228
rect 17727 7256 17739 7259
rect 20162 7256 20168 7268
rect 17727 7228 20168 7256
rect 17727 7225 17739 7228
rect 17681 7219 17739 7225
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 15160 7160 16773 7188
rect 15160 7148 15166 7160
rect 16761 7157 16773 7160
rect 16807 7188 16819 7191
rect 17543 7191 17601 7197
rect 17543 7188 17555 7191
rect 16807 7160 17555 7188
rect 16807 7157 16819 7160
rect 16761 7151 16819 7157
rect 17543 7157 17555 7160
rect 17589 7188 17601 7191
rect 18874 7188 18880 7200
rect 17589 7160 18880 7188
rect 17589 7157 17601 7160
rect 17543 7151 17601 7157
rect 18874 7148 18880 7160
rect 18932 7188 18938 7200
rect 20438 7188 20444 7200
rect 18932 7160 20444 7188
rect 18932 7148 18938 7160
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20625 7191 20683 7197
rect 20625 7157 20637 7191
rect 20671 7188 20683 7191
rect 20990 7188 20996 7200
rect 20671 7160 20996 7188
rect 20671 7157 20683 7160
rect 20625 7151 20683 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 1104 7098 26864 7120
rect 1104 7046 4169 7098
rect 4221 7046 4233 7098
rect 4285 7046 4297 7098
rect 4349 7046 4361 7098
rect 4413 7046 4425 7098
rect 4477 7046 10608 7098
rect 10660 7046 10672 7098
rect 10724 7046 10736 7098
rect 10788 7046 10800 7098
rect 10852 7046 10864 7098
rect 10916 7046 17047 7098
rect 17099 7046 17111 7098
rect 17163 7046 17175 7098
rect 17227 7046 17239 7098
rect 17291 7046 17303 7098
rect 17355 7046 23486 7098
rect 23538 7046 23550 7098
rect 23602 7046 23614 7098
rect 23666 7046 23678 7098
rect 23730 7046 23742 7098
rect 23794 7046 26864 7098
rect 1104 7024 26864 7046
rect 5261 6987 5319 6993
rect 5261 6953 5273 6987
rect 5307 6984 5319 6987
rect 5307 6956 5396 6984
rect 5307 6953 5319 6956
rect 5261 6947 5319 6953
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 3234 6848 3240 6860
rect 1627 6820 3240 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3375 6820 4077 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4706 6808 4712 6860
rect 4764 6808 4770 6860
rect 5368 6848 5396 6956
rect 5442 6944 5448 6996
rect 5500 6944 5506 6996
rect 8202 6944 8208 6996
rect 8260 6944 8266 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8352 6956 8677 6984
rect 8352 6944 8358 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8812 6956 9045 6984
rect 8812 6944 8818 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 9272 6956 9505 6984
rect 9272 6944 9278 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 5460 6916 5488 6944
rect 9508 6916 9536 6947
rect 10318 6944 10324 6996
rect 10376 6944 10382 6996
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10781 6987 10839 6993
rect 10781 6984 10793 6987
rect 10468 6956 10793 6984
rect 10468 6944 10474 6956
rect 10781 6953 10793 6956
rect 10827 6953 10839 6987
rect 10781 6947 10839 6953
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 11698 6984 11704 6996
rect 11655 6956 11704 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12032 6956 12357 6984
rect 12032 6944 12038 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 13630 6944 13636 6996
rect 13688 6944 13694 6996
rect 20530 6944 20536 6996
rect 20588 6944 20594 6996
rect 21450 6984 21456 6996
rect 20640 6956 21456 6984
rect 10229 6919 10287 6925
rect 5460 6888 5764 6916
rect 9508 6888 10180 6916
rect 5442 6848 5448 6860
rect 5368 6820 5448 6848
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 5736 6857 5764 6888
rect 5721 6851 5779 6857
rect 5500 6820 5672 6848
rect 5500 6808 5506 6820
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3050 6712 3056 6724
rect 2898 6684 3056 6712
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3620 6712 3648 6743
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3878 6780 3884 6792
rect 3752 6752 3884 6780
rect 3752 6740 3758 6752
rect 3878 6740 3884 6752
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4798 6780 4804 6792
rect 4295 6752 4804 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5258 6780 5264 6792
rect 5123 6752 5264 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5644 6789 5672 6820
rect 5721 6817 5733 6851
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5859 6820 6132 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 6104 6792 6132 6820
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 9180 6820 9229 6848
rect 9180 6808 9186 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9732 6820 9965 6848
rect 9732 6808 9738 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 4154 6712 4160 6724
rect 3620 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4341 6715 4399 6721
rect 4341 6681 4353 6715
rect 4387 6681 4399 6715
rect 4341 6675 4399 6681
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4356 6644 4384 6675
rect 4430 6672 4436 6724
rect 4488 6672 4494 6724
rect 4571 6715 4629 6721
rect 4571 6681 4583 6715
rect 4617 6712 4629 6715
rect 4706 6712 4712 6724
rect 4617 6684 4712 6712
rect 4617 6681 4629 6684
rect 4571 6675 4629 6681
rect 4706 6672 4712 6684
rect 4764 6712 4770 6724
rect 5445 6715 5503 6721
rect 5445 6712 5457 6715
rect 4764 6684 5457 6712
rect 4764 6672 4770 6684
rect 5445 6681 5457 6684
rect 5491 6681 5503 6715
rect 5644 6712 5672 6743
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8128 6712 8156 6743
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6782 9919 6783
rect 10045 6783 10103 6789
rect 9907 6754 9996 6782
rect 9907 6749 9919 6754
rect 9861 6743 9919 6749
rect 5644 6684 8156 6712
rect 9968 6712 9996 6754
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 10152 6780 10180 6888
rect 10229 6885 10241 6919
rect 10275 6916 10287 6919
rect 10594 6916 10600 6928
rect 10275 6888 10600 6916
rect 10275 6885 10287 6888
rect 10229 6879 10287 6885
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 10962 6916 10968 6928
rect 10704 6888 10968 6916
rect 10704 6848 10732 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11146 6876 11152 6928
rect 11204 6876 11210 6928
rect 11790 6916 11796 6928
rect 11256 6888 11796 6916
rect 10612 6820 10732 6848
rect 10091 6752 10180 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10612 6789 10640 6820
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 10284 6752 10517 6780
rect 10284 6740 10290 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11164 6789 11192 6876
rect 11256 6789 11284 6888
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 13596 6888 13676 6916
rect 13596 6876 13602 6888
rect 11606 6848 11612 6860
rect 11440 6820 11612 6848
rect 11440 6789 11468 6820
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 13648 6857 13676 6888
rect 20162 6876 20168 6928
rect 20220 6916 20226 6928
rect 20640 6916 20668 6956
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 20220 6888 20668 6916
rect 20220 6876 20226 6888
rect 13633 6851 13691 6857
rect 11808 6820 12572 6848
rect 11808 6789 11836 6820
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10744 6752 10885 6780
rect 10744 6740 10750 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12434 6780 12440 6792
rect 12115 6752 12440 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 9968 6684 10977 6712
rect 5445 6675 5503 6681
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 10965 6675 11023 6681
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4356 6616 4813 6644
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 5460 6644 5488 6675
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11532 6712 11560 6743
rect 12360 6721 12388 6752
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 12544 6721 12572 6820
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 16666 6848 16672 6860
rect 15887 6820 16672 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 19061 6851 19119 6857
rect 17460 6820 19012 6848
rect 17460 6808 17466 6820
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13136 6752 13553 6780
rect 13136 6740 13142 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13814 6740 13820 6792
rect 13872 6740 13878 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16298 6780 16304 6792
rect 16255 6752 16304 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 17678 6789 17684 6792
rect 17635 6783 17684 6789
rect 17635 6780 17647 6783
rect 17591 6752 17647 6780
rect 17635 6749 17647 6752
rect 17681 6749 17684 6783
rect 17635 6743 17684 6749
rect 17678 6740 17684 6743
rect 17736 6780 17742 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 17736 6752 18337 6780
rect 17736 6740 17742 6752
rect 18325 6749 18337 6752
rect 18371 6780 18383 6783
rect 18690 6780 18696 6792
rect 18371 6752 18696 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 18874 6740 18880 6792
rect 18932 6740 18938 6792
rect 18984 6780 19012 6820
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 19107 6820 20269 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 20257 6817 20269 6820
rect 20303 6848 20315 6851
rect 20303 6820 20760 6848
rect 20303 6817 20315 6820
rect 20257 6811 20315 6817
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 18984 6752 19257 6780
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 19978 6780 19984 6792
rect 19935 6752 19984 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6749 20683 6783
rect 20732 6780 20760 6820
rect 20990 6808 20996 6860
rect 21048 6808 21054 6860
rect 21450 6808 21456 6860
rect 21508 6848 21514 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21508 6820 22477 6848
rect 21508 6808 21514 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 21082 6780 21088 6792
rect 20732 6752 21088 6780
rect 20625 6743 20683 6749
rect 12329 6715 12388 6721
rect 11112 6684 12204 6712
rect 11112 6672 11118 6684
rect 5902 6644 5908 6656
rect 5460 6616 5908 6644
rect 4801 6607 4859 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 6052 6616 6101 6644
rect 6052 6604 6058 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 11974 6644 11980 6656
rect 8536 6616 11980 6644
rect 8536 6604 8542 6616
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12176 6653 12204 6684
rect 12329 6681 12341 6715
rect 12375 6684 12388 6715
rect 12529 6715 12587 6721
rect 12375 6681 12387 6684
rect 12329 6675 12387 6681
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 12986 6712 12992 6724
rect 12575 6684 12992 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 16942 6672 16948 6724
rect 17000 6672 17006 6724
rect 17402 6672 17408 6724
rect 17460 6712 17466 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 17460 6684 17785 6712
rect 17460 6672 17466 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 20640 6712 20668 6743
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 19208 6684 20668 6712
rect 19208 6672 19214 6684
rect 21910 6672 21916 6724
rect 21968 6672 21974 6724
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 13354 6604 13360 6656
rect 13412 6604 13418 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 19058 6644 19064 6656
rect 18104 6616 19064 6644
rect 18104 6604 18110 6616
rect 19058 6604 19064 6616
rect 19116 6644 19122 6656
rect 19978 6644 19984 6656
rect 19116 6616 19984 6644
rect 19116 6604 19122 6616
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 1104 6554 26864 6576
rect 1104 6502 4829 6554
rect 4881 6502 4893 6554
rect 4945 6502 4957 6554
rect 5009 6502 5021 6554
rect 5073 6502 5085 6554
rect 5137 6502 11268 6554
rect 11320 6502 11332 6554
rect 11384 6502 11396 6554
rect 11448 6502 11460 6554
rect 11512 6502 11524 6554
rect 11576 6502 17707 6554
rect 17759 6502 17771 6554
rect 17823 6502 17835 6554
rect 17887 6502 17899 6554
rect 17951 6502 17963 6554
rect 18015 6502 24146 6554
rect 24198 6502 24210 6554
rect 24262 6502 24274 6554
rect 24326 6502 24338 6554
rect 24390 6502 24402 6554
rect 24454 6502 26864 6554
rect 1104 6480 26864 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 4433 6443 4491 6449
rect 2455 6412 4384 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1596 6304 1624 6403
rect 3878 6372 3884 6384
rect 3450 6344 3884 6372
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 4356 6372 4384 6412
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4522 6440 4528 6452
rect 4479 6412 4528 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 5166 6440 5172 6452
rect 4856 6412 5172 6440
rect 4856 6400 4862 6412
rect 5166 6400 5172 6412
rect 5224 6440 5230 6452
rect 6086 6440 6092 6452
rect 5224 6412 6092 6440
rect 5224 6400 5230 6412
rect 6086 6400 6092 6412
rect 6144 6440 6150 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 6144 6412 7113 6440
rect 6144 6400 6150 6412
rect 7101 6409 7113 6412
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 9325 6443 9383 6449
rect 9325 6440 9337 6443
rect 8067 6412 9337 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 9325 6409 9337 6412
rect 9371 6440 9383 6443
rect 9490 6440 9496 6452
rect 9371 6412 9496 6440
rect 9371 6409 9383 6412
rect 9325 6403 9383 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10337 6443 10395 6449
rect 10337 6440 10349 6443
rect 10008 6412 10349 6440
rect 10008 6400 10014 6412
rect 10337 6409 10349 6412
rect 10383 6409 10395 6443
rect 10337 6403 10395 6409
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 10686 6400 10692 6452
rect 10744 6400 10750 6452
rect 16298 6400 16304 6452
rect 16356 6400 16362 6452
rect 16942 6400 16948 6452
rect 17000 6400 17006 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20128 6412 20637 6440
rect 20128 6400 20134 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 21910 6400 21916 6452
rect 21968 6400 21974 6452
rect 5442 6372 5448 6384
rect 4356 6344 5448 6372
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1596 6276 2145 6304
rect 1397 6267 1455 6273
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4798 6264 4804 6316
rect 4856 6264 4862 6316
rect 4908 6313 4936 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5537 6375 5595 6381
rect 5537 6341 5549 6375
rect 5583 6372 5595 6375
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 5583 6344 5825 6372
rect 5583 6341 5595 6344
rect 5537 6335 5595 6341
rect 5813 6341 5825 6344
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 5902 6332 5908 6384
rect 5960 6332 5966 6384
rect 7561 6375 7619 6381
rect 7561 6372 7573 6375
rect 6564 6344 7573 6372
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5258 6304 5264 6316
rect 5215 6276 5264 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 3786 6196 3792 6248
rect 3844 6236 3850 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3844 6208 3893 6236
rect 3844 6196 3850 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4488 6208 4721 6236
rect 4488 6196 4494 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 5092 6236 5120 6267
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5718 6304 5724 6316
rect 5675 6276 5724 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6564 6245 6592 6344
rect 7561 6341 7573 6344
rect 7607 6341 7619 6375
rect 7561 6335 7619 6341
rect 7653 6375 7711 6381
rect 7653 6341 7665 6375
rect 7699 6372 7711 6375
rect 8113 6375 8171 6381
rect 8113 6372 8125 6375
rect 7699 6344 8125 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 8113 6341 8125 6344
rect 8159 6372 8171 6375
rect 8202 6372 8208 6384
rect 8159 6344 8208 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 7282 6304 7288 6316
rect 6788 6276 7288 6304
rect 6788 6264 6794 6276
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7576 6304 7604 6335
rect 8202 6332 8208 6344
rect 8260 6372 8266 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 8260 6344 8585 6372
rect 8260 6332 8266 6344
rect 8573 6341 8585 6344
rect 8619 6341 8631 6375
rect 8573 6335 8631 6341
rect 9122 6332 9128 6384
rect 9180 6332 9186 6384
rect 9585 6375 9643 6381
rect 9585 6341 9597 6375
rect 9631 6372 9643 6375
rect 9674 6372 9680 6384
rect 9631 6344 9680 6372
rect 9631 6341 9643 6344
rect 9585 6335 9643 6341
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 10137 6375 10195 6381
rect 10137 6372 10149 6375
rect 9784 6344 10149 6372
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7576 6276 7849 6304
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7837 6267 7895 6273
rect 8036 6276 8309 6304
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5092 6208 6377 6236
rect 4709 6199 4767 6205
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 4724 6168 4752 6199
rect 5718 6168 5724 6180
rect 4724 6140 5724 6168
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6564 6168 6592 6199
rect 6638 6196 6644 6248
rect 6696 6196 6702 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 6914 6236 6920 6248
rect 6871 6208 6920 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 6914 6196 6920 6208
rect 6972 6236 6978 6248
rect 7466 6236 7472 6248
rect 6972 6208 7472 6236
rect 6972 6196 6978 6208
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8036 6168 8064 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8478 6264 8484 6316
rect 8536 6264 8542 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 6052 6140 6592 6168
rect 7300 6140 8064 6168
rect 6052 6128 6058 6140
rect 2222 6060 2228 6112
rect 2280 6060 2286 6112
rect 6178 6060 6184 6112
rect 6236 6060 6242 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7300 6109 7328 6140
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 6696 6072 7297 6100
rect 6696 6060 6702 6072
rect 7285 6069 7297 6072
rect 7331 6069 7343 6103
rect 7285 6063 7343 6069
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 8110 6100 8116 6112
rect 7524 6072 8116 6100
rect 7524 6060 7530 6072
rect 8110 6060 8116 6072
rect 8168 6100 8174 6112
rect 8772 6100 8800 6267
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9784 6304 9812 6344
rect 10137 6341 10149 6344
rect 10183 6341 10195 6375
rect 10612 6372 10640 6400
rect 17402 6372 17408 6384
rect 10612 6344 12434 6372
rect 10137 6335 10195 6341
rect 9692 6276 9812 6304
rect 9861 6310 9919 6313
rect 9861 6307 9996 6310
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9692 6236 9720 6276
rect 9861 6273 9873 6307
rect 9907 6304 9996 6307
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 9907 6282 10609 6304
rect 9907 6273 9919 6282
rect 9968 6276 10609 6282
rect 9861 6267 9919 6273
rect 9272 6208 9720 6236
rect 9272 6196 9278 6208
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 10134 6196 10140 6248
rect 10192 6236 10198 6248
rect 10410 6236 10416 6248
rect 10192 6208 10416 6236
rect 10192 6196 10198 6208
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10520 6177 10548 6276
rect 10597 6273 10609 6276
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 10505 6171 10563 6177
rect 9539 6140 10456 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 8168 6072 8800 6100
rect 9309 6103 9367 6109
rect 8168 6060 8174 6072
rect 9309 6069 9321 6103
rect 9355 6100 9367 6103
rect 9766 6100 9772 6112
rect 9355 6072 9772 6100
rect 9355 6069 9367 6072
rect 9309 6063 9367 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9876 6109 9904 6140
rect 9861 6103 9919 6109
rect 9861 6069 9873 6103
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 10045 6103 10103 6109
rect 10045 6069 10057 6103
rect 10091 6100 10103 6103
rect 10226 6100 10232 6112
rect 10091 6072 10232 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10318 6060 10324 6112
rect 10376 6060 10382 6112
rect 10428 6100 10456 6140
rect 10505 6137 10517 6171
rect 10551 6137 10563 6171
rect 10505 6131 10563 6137
rect 10796 6100 10824 6267
rect 12406 6168 12434 6344
rect 16408 6344 17408 6372
rect 15194 6264 15200 6316
rect 15252 6264 15258 6316
rect 16408 6313 16436 6344
rect 17402 6332 17408 6344
rect 17460 6332 17466 6384
rect 18874 6332 18880 6384
rect 18932 6372 18938 6384
rect 19889 6375 19947 6381
rect 18932 6344 19472 6372
rect 18932 6332 18938 6344
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6273 16451 6307
rect 16393 6267 16451 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 15212 6236 15240 6264
rect 15378 6236 15384 6248
rect 15212 6208 15384 6236
rect 15378 6196 15384 6208
rect 15436 6236 15442 6248
rect 17052 6236 17080 6267
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 19444 6313 19472 6344
rect 19889 6341 19901 6375
rect 19935 6372 19947 6375
rect 21082 6372 21088 6384
rect 19935 6344 21088 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 18748 6276 19257 6304
rect 18748 6264 18754 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 18322 6236 18328 6248
rect 15436 6208 18328 6236
rect 15436 6196 15442 6208
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 19337 6239 19395 6245
rect 19337 6205 19349 6239
rect 19383 6236 19395 6239
rect 19720 6236 19748 6267
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 20806 6304 20812 6316
rect 20036 6276 20812 6304
rect 20036 6264 20042 6276
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 21450 6304 21456 6316
rect 21315 6276 21456 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 21818 6264 21824 6316
rect 21876 6264 21882 6316
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 19383 6208 21189 6236
rect 19383 6205 19395 6208
rect 19337 6199 19395 6205
rect 21177 6205 21189 6208
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 20714 6168 20720 6180
rect 12406 6140 20720 6168
rect 20714 6128 20720 6140
rect 20772 6128 20778 6180
rect 20898 6128 20904 6180
rect 20956 6128 20962 6180
rect 10428 6072 10824 6100
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 15068 6072 15117 6100
rect 15068 6060 15074 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 19521 6103 19579 6109
rect 19521 6069 19533 6103
rect 19567 6100 19579 6103
rect 19610 6100 19616 6112
rect 19567 6072 19616 6100
rect 19567 6069 19579 6072
rect 19521 6063 19579 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 1104 6010 26864 6032
rect 1104 5958 4169 6010
rect 4221 5958 4233 6010
rect 4285 5958 4297 6010
rect 4349 5958 4361 6010
rect 4413 5958 4425 6010
rect 4477 5958 10608 6010
rect 10660 5958 10672 6010
rect 10724 5958 10736 6010
rect 10788 5958 10800 6010
rect 10852 5958 10864 6010
rect 10916 5958 17047 6010
rect 17099 5958 17111 6010
rect 17163 5958 17175 6010
rect 17227 5958 17239 6010
rect 17291 5958 17303 6010
rect 17355 5958 23486 6010
rect 23538 5958 23550 6010
rect 23602 5958 23614 6010
rect 23666 5958 23678 6010
rect 23730 5958 23742 6010
rect 23794 5958 26864 6010
rect 1104 5936 26864 5958
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 4672 5868 5181 5896
rect 4672 5856 4678 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 5169 5859 5227 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 5316 5868 5549 5896
rect 5316 5856 5322 5868
rect 5537 5865 5549 5868
rect 5583 5865 5595 5899
rect 5537 5859 5595 5865
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6270 5896 6276 5908
rect 6227 5868 6276 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 9674 5856 9680 5908
rect 9732 5856 9738 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 12894 5896 12900 5908
rect 10376 5868 12900 5896
rect 10376 5856 10382 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 25685 5899 25743 5905
rect 25685 5896 25697 5899
rect 13044 5868 25697 5896
rect 13044 5856 13050 5868
rect 25685 5865 25697 5868
rect 25731 5865 25743 5899
rect 25685 5859 25743 5865
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5797 5043 5831
rect 4985 5791 5043 5797
rect 6411 5831 6469 5837
rect 6411 5797 6423 5831
rect 6457 5828 6469 5831
rect 6546 5828 6552 5840
rect 6457 5800 6552 5828
rect 6457 5797 6469 5800
rect 6411 5791 6469 5797
rect 5000 5760 5028 5791
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 9585 5831 9643 5837
rect 9585 5797 9597 5831
rect 9631 5828 9643 5831
rect 9858 5828 9864 5840
rect 9631 5800 9864 5828
rect 9631 5797 9643 5800
rect 9585 5791 9643 5797
rect 9858 5788 9864 5800
rect 9916 5828 9922 5840
rect 10152 5828 10180 5856
rect 9916 5800 10180 5828
rect 9916 5788 9922 5800
rect 5166 5760 5172 5772
rect 5000 5732 5172 5760
rect 5166 5720 5172 5732
rect 5224 5760 5230 5772
rect 5350 5760 5356 5772
rect 5224 5732 5356 5760
rect 5224 5720 5230 5732
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 6914 5760 6920 5772
rect 6104 5732 6920 5760
rect 5626 5692 5632 5704
rect 5276 5664 5632 5692
rect 2222 5584 2228 5636
rect 2280 5624 2286 5636
rect 5153 5627 5211 5633
rect 2280 5596 2774 5624
rect 2280 5584 2286 5596
rect 2746 5556 2774 5596
rect 5153 5593 5165 5627
rect 5199 5624 5211 5627
rect 5276 5624 5304 5664
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6104 5701 6132 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 10336 5760 10364 5856
rect 13906 5788 13912 5840
rect 13964 5828 13970 5840
rect 14139 5831 14197 5837
rect 14139 5828 14151 5831
rect 13964 5800 14151 5828
rect 13964 5788 13970 5800
rect 14139 5797 14151 5800
rect 14185 5797 14197 5831
rect 14139 5791 14197 5797
rect 19334 5788 19340 5840
rect 19392 5788 19398 5840
rect 20070 5828 20076 5840
rect 19444 5800 20076 5828
rect 9416 5732 10364 5760
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6730 5692 6736 5704
rect 6595 5664 6736 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 5199 5596 5304 5624
rect 5353 5627 5411 5633
rect 5199 5593 5211 5596
rect 5153 5587 5211 5593
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5442 5624 5448 5636
rect 5399 5596 5448 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 6288 5624 6316 5655
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9416 5701 9444 5732
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 8996 5664 9321 5692
rect 8996 5652 9002 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9548 5664 9965 5692
rect 9548 5652 9554 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16666 5692 16672 5704
rect 15979 5664 16672 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16666 5652 16672 5664
rect 16724 5692 16730 5704
rect 19337 5695 19395 5701
rect 16724 5664 17816 5692
rect 16724 5652 16730 5664
rect 6052 5596 6316 5624
rect 6052 5584 6058 5596
rect 9214 5584 9220 5636
rect 9272 5624 9278 5636
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 9272 5596 9597 5624
rect 9272 5584 9278 5596
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 9677 5627 9735 5633
rect 9677 5593 9689 5627
rect 9723 5593 9735 5627
rect 9677 5587 9735 5593
rect 7190 5556 7196 5568
rect 2746 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9692 5556 9720 5587
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 9824 5596 9873 5624
rect 9824 5584 9830 5596
rect 9861 5593 9873 5596
rect 9907 5624 9919 5627
rect 13354 5624 13360 5636
rect 9907 5596 13360 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 15010 5584 15016 5636
rect 15068 5584 15074 5636
rect 17788 5633 17816 5664
rect 19337 5661 19349 5695
rect 19383 5692 19395 5695
rect 19444 5692 19472 5800
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 20346 5760 20352 5772
rect 19720 5732 20352 5760
rect 19383 5664 19472 5692
rect 19383 5661 19395 5664
rect 19337 5655 19395 5661
rect 19518 5652 19524 5704
rect 19576 5652 19582 5704
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 19720 5701 19748 5732
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 25777 5695 25835 5701
rect 25777 5661 25789 5695
rect 25823 5692 25835 5695
rect 26326 5692 26332 5704
rect 25823 5664 26332 5692
rect 25823 5661 25835 5664
rect 25777 5655 25835 5661
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5593 16083 5627
rect 16025 5587 16083 5593
rect 17773 5627 17831 5633
rect 17773 5593 17785 5627
rect 17819 5624 17831 5627
rect 19150 5624 19156 5636
rect 17819 5596 19156 5624
rect 17819 5593 17831 5596
rect 17773 5587 17831 5593
rect 9548 5528 9720 5556
rect 9548 5516 9554 5528
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 16040 5556 16068 5587
rect 19150 5584 19156 5596
rect 19208 5584 19214 5636
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19797 5627 19855 5633
rect 19797 5624 19809 5627
rect 19484 5596 19809 5624
rect 19484 5584 19490 5596
rect 19797 5593 19809 5596
rect 19843 5593 19855 5627
rect 19797 5587 19855 5593
rect 18230 5556 18236 5568
rect 14424 5528 18236 5556
rect 14424 5516 14430 5528
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 19904 5556 19932 5655
rect 26326 5652 26332 5664
rect 26384 5652 26390 5704
rect 19576 5528 19932 5556
rect 19576 5516 19582 5528
rect 1104 5466 26864 5488
rect 1104 5414 4829 5466
rect 4881 5414 4893 5466
rect 4945 5414 4957 5466
rect 5009 5414 5021 5466
rect 5073 5414 5085 5466
rect 5137 5414 11268 5466
rect 11320 5414 11332 5466
rect 11384 5414 11396 5466
rect 11448 5414 11460 5466
rect 11512 5414 11524 5466
rect 11576 5414 17707 5466
rect 17759 5414 17771 5466
rect 17823 5414 17835 5466
rect 17887 5414 17899 5466
rect 17951 5414 17963 5466
rect 18015 5414 24146 5466
rect 24198 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 26864 5466
rect 1104 5392 26864 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 5981 5355 6039 5361
rect 5981 5321 5993 5355
rect 6027 5352 6039 5355
rect 6270 5352 6276 5364
rect 6027 5324 6276 5352
rect 6027 5321 6039 5324
rect 5981 5315 6039 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 14277 5355 14335 5361
rect 13556 5324 13860 5352
rect 6181 5287 6239 5293
rect 6181 5253 6193 5287
rect 6227 5284 6239 5287
rect 6914 5284 6920 5296
rect 6227 5256 6920 5284
rect 6227 5253 6239 5256
rect 6181 5247 6239 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 9582 5244 9588 5296
rect 9640 5244 9646 5296
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 1636 5188 2145 5216
rect 1636 5176 1642 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 9122 5216 9128 5228
rect 2547 5188 9128 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 9122 5176 9128 5188
rect 9180 5216 9186 5228
rect 9490 5216 9496 5228
rect 9180 5188 9496 5216
rect 9180 5176 9186 5188
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 12434 5176 12440 5228
rect 12492 5176 12498 5228
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13136 5188 13277 5216
rect 13136 5176 13142 5188
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 13446 5176 13452 5228
rect 13504 5216 13510 5228
rect 13556 5225 13584 5324
rect 13630 5244 13636 5296
rect 13688 5244 13694 5296
rect 13832 5284 13860 5324
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14323 5324 15332 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 13832 5256 14780 5284
rect 13832 5225 13860 5256
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13504 5188 13553 5216
rect 13504 5176 13510 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13725 5219 13783 5225
rect 13725 5206 13737 5219
rect 13541 5179 13599 5185
rect 13648 5185 13737 5206
rect 13771 5185 13783 5219
rect 13648 5179 13783 5185
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 13648 5178 13768 5179
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5148 2283 5151
rect 9214 5148 9220 5160
rect 2271 5120 9220 5148
rect 2271 5117 2283 5120
rect 2225 5111 2283 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 13648 5148 13676 5178
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 14056 5188 14105 5216
rect 14056 5176 14062 5188
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 14139 5188 14657 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14752 5216 14780 5256
rect 14752 5188 14872 5216
rect 14645 5179 14703 5185
rect 13906 5148 13912 5160
rect 13648 5120 13912 5148
rect 13906 5108 13912 5120
rect 13964 5148 13970 5160
rect 14844 5157 14872 5188
rect 15102 5176 15108 5228
rect 15160 5176 15166 5228
rect 15304 5225 15332 5324
rect 19334 5312 19340 5364
rect 19392 5312 19398 5364
rect 19153 5287 19211 5293
rect 19153 5253 19165 5287
rect 19199 5284 19211 5287
rect 19352 5284 19380 5312
rect 19199 5256 19380 5284
rect 19199 5253 19211 5256
rect 19153 5247 19211 5253
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 16574 5216 16580 5228
rect 15335 5188 16580 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 19334 5176 19340 5228
rect 19392 5176 19398 5228
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 19610 5216 19616 5228
rect 19475 5188 19616 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 13964 5120 14565 5148
rect 13964 5108 13970 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 12158 5040 12164 5092
rect 12216 5080 12222 5092
rect 13262 5080 13268 5092
rect 12216 5052 13268 5080
rect 12216 5040 12222 5052
rect 13262 5040 13268 5052
rect 13320 5080 13326 5092
rect 13403 5083 13461 5089
rect 13403 5080 13415 5083
rect 13320 5052 13415 5080
rect 13320 5040 13326 5052
rect 13403 5049 13415 5052
rect 13449 5080 13461 5083
rect 14752 5080 14780 5111
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 19904 5148 19932 5179
rect 20898 5148 20904 5160
rect 18380 5120 20904 5148
rect 18380 5108 18386 5120
rect 20898 5108 20904 5120
rect 20956 5148 20962 5160
rect 21818 5148 21824 5160
rect 20956 5120 21824 5148
rect 20956 5108 20962 5120
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 13449 5052 14780 5080
rect 13449 5049 13461 5052
rect 13403 5043 13461 5049
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 8294 4972 8300 5024
rect 8352 4972 8358 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 10560 4984 12633 5012
rect 10560 4972 10566 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 13078 4972 13084 5024
rect 13136 5012 13142 5024
rect 13998 5012 14004 5024
rect 13136 4984 14004 5012
rect 13136 4972 13142 4984
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14108 5021 14136 5052
rect 14093 5015 14151 5021
rect 14093 4981 14105 5015
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 15010 4972 15016 5024
rect 15068 4972 15074 5024
rect 15102 4972 15108 5024
rect 15160 5012 15166 5024
rect 15197 5015 15255 5021
rect 15197 5012 15209 5015
rect 15160 4984 15209 5012
rect 15160 4972 15166 4984
rect 15197 4981 15209 4984
rect 15243 4981 15255 5015
rect 15197 4975 15255 4981
rect 19153 5015 19211 5021
rect 19153 4981 19165 5015
rect 19199 5012 19211 5015
rect 19242 5012 19248 5024
rect 19199 4984 19248 5012
rect 19199 4981 19211 4984
rect 19153 4975 19211 4981
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 19978 4972 19984 5024
rect 20036 4972 20042 5024
rect 1104 4922 26864 4944
rect 1104 4870 4169 4922
rect 4221 4870 4233 4922
rect 4285 4870 4297 4922
rect 4349 4870 4361 4922
rect 4413 4870 4425 4922
rect 4477 4870 10608 4922
rect 10660 4870 10672 4922
rect 10724 4870 10736 4922
rect 10788 4870 10800 4922
rect 10852 4870 10864 4922
rect 10916 4870 17047 4922
rect 17099 4870 17111 4922
rect 17163 4870 17175 4922
rect 17227 4870 17239 4922
rect 17291 4870 17303 4922
rect 17355 4870 23486 4922
rect 23538 4870 23550 4922
rect 23602 4870 23614 4922
rect 23666 4870 23678 4922
rect 23730 4870 23742 4922
rect 23794 4870 26864 4922
rect 1104 4848 26864 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 8110 4768 8116 4820
rect 8168 4768 8174 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 11054 4808 11060 4820
rect 10100 4780 11060 4808
rect 10100 4768 10106 4780
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 12728 4780 13492 4808
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6236 4644 6653 4672
rect 6236 4632 6242 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 8352 4644 10149 4672
rect 8352 4632 8358 4644
rect 10137 4641 10149 4644
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 10502 4632 10508 4684
rect 10560 4632 10566 4684
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4764 4576 4813 4604
rect 4764 4564 4770 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 5166 4604 5172 4616
rect 5031 4576 5172 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8386 4604 8392 4616
rect 8076 4576 8392 4604
rect 8076 4564 8082 4576
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 12728 4613 12756 4780
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 13136 4712 13400 4740
rect 13136 4700 13142 4712
rect 13004 4644 13308 4672
rect 13004 4613 13032 4644
rect 13280 4616 13308 4644
rect 11931 4607 11989 4613
rect 11931 4573 11943 4607
rect 11977 4604 11989 4607
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 11977 4576 12725 4604
rect 11977 4573 11989 4576
rect 11931 4567 11989 4573
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 13078 4564 13084 4616
rect 13136 4564 13142 4616
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 13372 4604 13400 4712
rect 13464 4672 13492 4780
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13596 4780 13737 4808
rect 13596 4768 13602 4780
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 13725 4771 13783 4777
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 15562 4808 15568 4820
rect 14691 4780 15568 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 16485 4811 16543 4817
rect 16485 4777 16497 4811
rect 16531 4808 16543 4811
rect 17402 4808 17408 4820
rect 16531 4780 17408 4808
rect 16531 4777 16543 4780
rect 16485 4771 16543 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 21039 4811 21097 4817
rect 21039 4808 21051 4811
rect 20864 4780 21051 4808
rect 20864 4768 20870 4780
rect 21039 4777 21051 4780
rect 21085 4777 21097 4811
rect 21039 4771 21097 4777
rect 18230 4740 18236 4752
rect 14200 4712 16988 4740
rect 14200 4672 14228 4712
rect 14737 4675 14795 4681
rect 14737 4672 14749 4675
rect 13464 4644 14228 4672
rect 14292 4644 14749 4672
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 13372 4576 13461 4604
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 13906 4564 13912 4616
rect 13964 4564 13970 4616
rect 14090 4564 14096 4616
rect 14148 4564 14154 4616
rect 14292 4613 14320 4644
rect 14737 4641 14749 4644
rect 14783 4641 14795 4675
rect 15102 4672 15108 4684
rect 14737 4635 14795 4641
rect 14844 4644 15108 4672
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14844 4604 14872 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4672 16359 4675
rect 16574 4672 16580 4684
rect 16347 4644 16580 4672
rect 16347 4641 16359 4644
rect 16301 4635 16359 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 16960 4681 16988 4712
rect 17052 4712 18236 4740
rect 17052 4684 17080 4712
rect 18230 4700 18236 4712
rect 18288 4700 18294 4752
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 16945 4635 17003 4641
rect 14507 4576 14872 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14918 4564 14924 4616
rect 14976 4564 14982 4616
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 15068 4576 15209 4604
rect 15068 4564 15074 4576
rect 15197 4573 15209 4576
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 4430 4496 4436 4548
rect 4488 4536 4494 4548
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4488 4508 5365 4536
rect 4488 4496 4494 4508
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 5353 4499 5411 4505
rect 5534 4496 5540 4548
rect 5592 4496 5598 4548
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4536 5779 4539
rect 6270 4536 6276 4548
rect 5767 4508 6276 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 6270 4496 6276 4508
rect 6328 4496 6334 4548
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 7866 4508 8309 4536
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 12805 4539 12863 4545
rect 8297 4499 8355 4505
rect 10796 4508 10902 4536
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 4522 4468 4528 4480
rect 4304 4440 4528 4468
rect 4304 4428 4310 4440
rect 4522 4428 4528 4440
rect 4580 4468 4586 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4580 4440 4905 4468
rect 4580 4428 4586 4440
rect 4893 4437 4905 4440
rect 4939 4437 4951 4471
rect 4893 4431 4951 4437
rect 9950 4428 9956 4480
rect 10008 4428 10014 4480
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10796 4468 10824 4508
rect 12805 4505 12817 4539
rect 12851 4536 12863 4539
rect 12894 4536 12900 4548
rect 12851 4508 12900 4536
rect 12851 4505 12863 4508
rect 12805 4499 12863 4505
rect 12894 4496 12900 4508
rect 12952 4536 12958 4548
rect 13541 4539 13599 4545
rect 12952 4508 13492 4536
rect 12952 4496 12958 4508
rect 10284 4440 10824 4468
rect 10284 4428 10290 4440
rect 12526 4428 12532 4480
rect 12584 4428 12590 4480
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13044 4440 13369 4468
rect 13044 4428 13050 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13464 4468 13492 4508
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 13924 4536 13952 4564
rect 13587 4508 13952 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 14366 4496 14372 4548
rect 14424 4496 14430 4548
rect 15856 4536 15884 4567
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16758 4604 16764 4616
rect 16264 4576 16764 4604
rect 16264 4564 16270 4576
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16960 4604 16988 4635
rect 17034 4632 17040 4684
rect 17092 4632 17098 4684
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 18046 4672 18052 4684
rect 17175 4644 18052 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 19150 4632 19156 4684
rect 19208 4672 19214 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 19208 4644 19257 4672
rect 19208 4632 19214 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19484 4644 19625 4672
rect 19484 4632 19490 4644
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16960 4576 17509 4604
rect 16853 4567 16911 4573
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 18414 4604 18420 4616
rect 17543 4576 18420 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 16868 4536 16896 4567
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 18049 4539 18107 4545
rect 18049 4536 18061 4539
rect 15028 4508 18061 4536
rect 13741 4471 13799 4477
rect 13741 4468 13753 4471
rect 13464 4440 13753 4468
rect 13357 4431 13415 4437
rect 13741 4437 13753 4440
rect 13787 4437 13799 4471
rect 13741 4431 13799 4437
rect 13906 4428 13912 4480
rect 13964 4468 13970 4480
rect 15028 4468 15056 4508
rect 18049 4505 18061 4508
rect 18095 4505 18107 4539
rect 18049 4499 18107 4505
rect 18230 4496 18236 4548
rect 18288 4496 18294 4548
rect 19978 4496 19984 4548
rect 20036 4496 20042 4548
rect 13964 4440 15056 4468
rect 15105 4471 15163 4477
rect 13964 4428 13970 4440
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 15654 4468 15660 4480
rect 15151 4440 15660 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 15654 4428 15660 4440
rect 15712 4468 15718 4480
rect 15749 4471 15807 4477
rect 15749 4468 15761 4471
rect 15712 4440 15761 4468
rect 15712 4428 15718 4440
rect 15749 4437 15761 4440
rect 15795 4437 15807 4471
rect 15749 4431 15807 4437
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16942 4468 16948 4480
rect 16715 4440 16948 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17218 4428 17224 4480
rect 17276 4468 17282 4480
rect 17405 4471 17463 4477
rect 17405 4468 17417 4471
rect 17276 4440 17417 4468
rect 17276 4428 17282 4440
rect 17405 4437 17417 4440
rect 17451 4437 17463 4471
rect 17405 4431 17463 4437
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 18196 4440 18429 4468
rect 18196 4428 18202 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 1104 4378 26864 4400
rect 1104 4326 4829 4378
rect 4881 4326 4893 4378
rect 4945 4326 4957 4378
rect 5009 4326 5021 4378
rect 5073 4326 5085 4378
rect 5137 4326 11268 4378
rect 11320 4326 11332 4378
rect 11384 4326 11396 4378
rect 11448 4326 11460 4378
rect 11512 4326 11524 4378
rect 11576 4326 17707 4378
rect 17759 4326 17771 4378
rect 17823 4326 17835 4378
rect 17887 4326 17899 4378
rect 17951 4326 17963 4378
rect 18015 4326 24146 4378
rect 24198 4326 24210 4378
rect 24262 4326 24274 4378
rect 24326 4326 24338 4378
rect 24390 4326 24402 4378
rect 24454 4326 26864 4378
rect 1104 4304 26864 4326
rect 4246 4224 4252 4276
rect 4304 4224 4310 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10100 4236 10609 4264
rect 10100 4224 10106 4236
rect 10597 4233 10609 4236
rect 10643 4233 10655 4267
rect 11970 4267 12028 4273
rect 11970 4264 11982 4267
rect 10597 4227 10655 4233
rect 11164 4236 11982 4264
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 4154 4196 4160 4208
rect 4111 4168 4160 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 4709 4199 4767 4205
rect 4264 4168 4660 4196
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 4264 4128 4292 4168
rect 3752 4100 4292 4128
rect 4341 4131 4399 4137
rect 3752 4088 3758 4100
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 4430 4128 4436 4140
rect 4387 4100 4436 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4632 4128 4660 4168
rect 4709 4165 4721 4199
rect 4755 4196 4767 4199
rect 5077 4199 5135 4205
rect 5077 4196 5089 4199
rect 4755 4168 5089 4196
rect 4755 4165 4767 4168
rect 4709 4159 4767 4165
rect 5077 4165 5089 4168
rect 5123 4165 5135 4199
rect 5077 4159 5135 4165
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5997 4199 6055 4205
rect 5997 4196 6009 4199
rect 5224 4168 6009 4196
rect 5224 4156 5230 4168
rect 5997 4165 6009 4168
rect 6043 4165 6055 4199
rect 5997 4159 6055 4165
rect 6362 4156 6368 4208
rect 6420 4196 6426 4208
rect 8294 4196 8300 4208
rect 6420 4168 6868 4196
rect 6420 4156 6426 4168
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4632 4100 4997 4128
rect 4525 4091 4583 4097
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5031 4100 5672 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 4540 4060 4568 4091
rect 4706 4060 4712 4072
rect 4540 4032 4712 4060
rect 4706 4020 4712 4032
rect 4764 4060 4770 4072
rect 5644 4060 5672 4100
rect 5718 4088 5724 4140
rect 5776 4088 5782 4140
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6730 4088 6736 4140
rect 6788 4088 6794 4140
rect 6840 4128 6868 4168
rect 8128 4168 8300 4196
rect 8128 4137 8156 4168
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 8846 4156 8852 4208
rect 8904 4156 8910 4208
rect 10229 4199 10287 4205
rect 10229 4165 10241 4199
rect 10275 4196 10287 4199
rect 11164 4196 11192 4236
rect 11970 4233 11982 4236
rect 12016 4233 12028 4267
rect 12526 4264 12532 4276
rect 11970 4227 12028 4233
rect 12084 4236 12532 4264
rect 12084 4205 12112 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 12676 4236 13492 4264
rect 12676 4224 12682 4236
rect 12069 4199 12127 4205
rect 10275 4168 11192 4196
rect 11440 4168 11652 4196
rect 10275 4165 10287 4168
rect 10229 4159 10287 4165
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 6840 4100 8125 4128
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 10410 4088 10416 4140
rect 10468 4088 10474 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11440 4128 11468 4168
rect 10551 4100 11468 4128
rect 11517 4131 11575 4137
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 11517 4097 11529 4131
rect 11563 4097 11575 4131
rect 11624 4128 11652 4168
rect 12069 4165 12081 4199
rect 12115 4165 12127 4199
rect 12069 4159 12127 4165
rect 12345 4199 12403 4205
rect 12345 4165 12357 4199
rect 12391 4196 12403 4199
rect 12986 4196 12992 4208
rect 12391 4168 12992 4196
rect 12391 4165 12403 4168
rect 12345 4159 12403 4165
rect 12986 4156 12992 4168
rect 13044 4156 13050 4208
rect 13354 4196 13360 4208
rect 13096 4168 13360 4196
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11624 4100 11805 4128
rect 11517 4091 11575 4097
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12434 4128 12440 4140
rect 11931 4100 12440 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 8018 4060 8024 4072
rect 4764 4032 5028 4060
rect 5644 4032 8024 4060
rect 4764 4020 4770 4032
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 4893 3995 4951 4001
rect 4893 3992 4905 3995
rect 4672 3964 4905 3992
rect 4672 3952 4678 3964
rect 4893 3961 4905 3964
rect 4939 3961 4951 3995
rect 5000 3992 5028 4032
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8478 4060 8484 4072
rect 8435 4032 8484 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9824 4032 10149 4060
rect 9824 4020 9830 4032
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 11112 4032 11161 4060
rect 11112 4020 11118 4032
rect 11149 4029 11161 4032
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 6638 3992 6644 4004
rect 5000 3964 6644 3992
rect 4893 3955 4951 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 11532 3992 11560 4091
rect 11808 4060 11836 4091
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11808 4032 12173 4060
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 9640 3964 11560 3992
rect 12452 3992 12480 4088
rect 12544 4060 12572 4091
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12805 4131 12863 4137
rect 12805 4128 12817 4131
rect 12768 4100 12817 4128
rect 12768 4088 12774 4100
rect 12805 4097 12817 4100
rect 12851 4128 12863 4131
rect 13096 4128 13124 4168
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 13464 4205 13492 4236
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14987 4267 15045 4273
rect 14987 4264 14999 4267
rect 13964 4236 14999 4264
rect 13964 4224 13970 4236
rect 14987 4233 14999 4236
rect 15033 4233 15045 4267
rect 14987 4227 15045 4233
rect 15120 4236 17816 4264
rect 13449 4199 13507 4205
rect 13449 4165 13461 4199
rect 13495 4165 13507 4199
rect 13449 4159 13507 4165
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 12851 4100 13124 4128
rect 13188 4100 13277 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 12894 4060 12900 4072
rect 12544 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 13188 4069 13216 4100
rect 13265 4097 13277 4100
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4029 13231 4063
rect 13464 4060 13492 4159
rect 14090 4156 14096 4208
rect 14148 4196 14154 4208
rect 15120 4196 15148 4236
rect 14148 4168 15148 4196
rect 15197 4199 15255 4205
rect 14148 4156 14154 4168
rect 15197 4165 15209 4199
rect 15243 4196 15255 4199
rect 15470 4196 15476 4208
rect 15243 4168 15476 4196
rect 15243 4165 15255 4168
rect 15197 4159 15255 4165
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 16206 4196 16212 4208
rect 15580 4168 16212 4196
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 15028 4100 15301 4128
rect 14918 4060 14924 4072
rect 13464 4032 14924 4060
rect 13173 4023 13231 4029
rect 13446 3992 13452 4004
rect 12452 3964 13452 3992
rect 9640 3952 9646 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 14844 4001 14872 4032
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 14829 3995 14887 4001
rect 14829 3961 14841 3995
rect 14875 3961 14887 3995
rect 14829 3955 14887 3961
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 4028 3896 4077 3924
rect 4028 3884 4034 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4212 3896 4721 3924
rect 4212 3884 4218 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 6178 3884 6184 3936
rect 6236 3884 6242 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 9766 3924 9772 3936
rect 6788 3896 9772 3924
rect 6788 3884 6794 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 10410 3924 10416 3936
rect 10275 3896 10416 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 11606 3884 11612 3936
rect 11664 3884 11670 3936
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13412 3896 13645 3924
rect 13412 3884 13418 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 15028 3933 15056 4100
rect 15289 4097 15301 4100
rect 15335 4128 15347 4131
rect 15580 4128 15608 4168
rect 16206 4156 16212 4168
rect 16264 4156 16270 4208
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 17680 4199 17738 4205
rect 16816 4168 17586 4196
rect 16816 4156 16822 4168
rect 15335 4100 15608 4128
rect 15335 4097 15347 4100
rect 15289 4091 15347 4097
rect 15654 4088 15660 4140
rect 15712 4088 15718 4140
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 16960 4060 16988 4091
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 17218 4088 17224 4140
rect 17276 4088 17282 4140
rect 17558 4137 17586 4168
rect 17680 4165 17692 4199
rect 17726 4196 17738 4199
rect 17788 4196 17816 4236
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 18141 4267 18199 4273
rect 18141 4264 18153 4267
rect 18104 4236 18153 4264
rect 18104 4224 18110 4236
rect 18141 4233 18153 4236
rect 18187 4233 18199 4267
rect 18141 4227 18199 4233
rect 20438 4224 20444 4276
rect 20496 4264 20502 4276
rect 20579 4267 20637 4273
rect 20579 4264 20591 4267
rect 20496 4236 20591 4264
rect 20496 4224 20502 4236
rect 20579 4233 20591 4236
rect 20625 4233 20637 4267
rect 20579 4227 20637 4233
rect 20809 4199 20867 4205
rect 20809 4196 20821 4199
rect 17726 4168 17816 4196
rect 20194 4168 20821 4196
rect 17726 4165 17738 4168
rect 17680 4159 17738 4165
rect 20809 4165 20821 4168
rect 20855 4165 20867 4199
rect 20809 4159 20867 4165
rect 17558 4131 17621 4137
rect 17558 4098 17575 4131
rect 17563 4097 17575 4098
rect 17609 4128 17621 4131
rect 17609 4098 17632 4128
rect 17609 4097 17621 4098
rect 17563 4091 17621 4097
rect 17770 4088 17776 4140
rect 17828 4088 17834 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18138 4128 18144 4140
rect 17911 4100 18144 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 18288 4100 18337 4128
rect 18288 4088 18294 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 18414 4088 18420 4140
rect 18472 4088 18478 4140
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 19058 4128 19064 4140
rect 18831 4100 19064 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 17310 4060 17316 4072
rect 16500 4032 17316 4060
rect 15841 3995 15899 4001
rect 15841 3961 15853 3995
rect 15887 3992 15899 3995
rect 16114 3992 16120 4004
rect 15887 3964 16120 3992
rect 15887 3961 15899 3964
rect 15841 3955 15899 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14792 3896 15025 3924
rect 14792 3884 14798 3896
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 16500 3924 16528 4032
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 17402 4020 17408 4072
rect 17460 4020 17466 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 17512 4032 18521 4060
rect 16574 3952 16580 4004
rect 16632 3992 16638 4004
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 16632 3964 17141 3992
rect 16632 3952 16638 3964
rect 17129 3961 17141 3964
rect 17175 3992 17187 3995
rect 17512 3992 17540 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 18414 3992 18420 4004
rect 17175 3964 17540 3992
rect 17604 3964 18420 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 15528 3896 16528 3924
rect 15528 3884 15534 3896
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17604 3924 17632 3964
rect 18414 3952 18420 3964
rect 18472 3992 18478 4004
rect 18616 3992 18644 4091
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19242 4128 19248 4140
rect 19199 4100 19248 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 18472 3964 18644 3992
rect 18472 3952 18478 3964
rect 26326 3952 26332 4004
rect 26384 3952 26390 4004
rect 17368 3896 17632 3924
rect 17368 3884 17374 3896
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17736 3896 18061 3924
rect 17736 3884 17742 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 1104 3834 26864 3856
rect 1104 3782 4169 3834
rect 4221 3782 4233 3834
rect 4285 3782 4297 3834
rect 4349 3782 4361 3834
rect 4413 3782 4425 3834
rect 4477 3782 10608 3834
rect 10660 3782 10672 3834
rect 10724 3782 10736 3834
rect 10788 3782 10800 3834
rect 10852 3782 10864 3834
rect 10916 3782 17047 3834
rect 17099 3782 17111 3834
rect 17163 3782 17175 3834
rect 17227 3782 17239 3834
rect 17291 3782 17303 3834
rect 17355 3782 23486 3834
rect 23538 3782 23550 3834
rect 23602 3782 23614 3834
rect 23666 3782 23678 3834
rect 23730 3782 23742 3834
rect 23794 3782 26864 3834
rect 1104 3760 26864 3782
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5718 3720 5724 3732
rect 5583 3692 5724 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 9033 3723 9091 3729
rect 9033 3689 9045 3723
rect 9079 3720 9091 3723
rect 10226 3720 10232 3732
rect 9079 3692 10232 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 11839 3723 11897 3729
rect 11839 3689 11851 3723
rect 11885 3720 11897 3723
rect 12158 3720 12164 3732
rect 11885 3692 12164 3720
rect 11885 3689 11897 3692
rect 11839 3683 11897 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 13596 3692 14197 3720
rect 13596 3680 13602 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 13725 3655 13783 3661
rect 13725 3621 13737 3655
rect 13771 3621 13783 3655
rect 13725 3615 13783 3621
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 4062 3584 4068 3596
rect 3835 3556 4068 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 6362 3584 6368 3596
rect 4120 3556 6368 3584
rect 4120 3544 4126 3556
rect 6362 3544 6368 3556
rect 6420 3584 6426 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6420 3556 6745 3584
rect 6420 3544 6426 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 8352 3556 10057 3584
rect 8352 3544 8358 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 12986 3584 12992 3596
rect 12851 3556 12992 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13740 3584 13768 3615
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 13127 3556 13584 3584
rect 13740 3556 15577 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3694 3516 3700 3528
rect 3467 3488 3700 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4246 3516 4252 3528
rect 4203 3488 4252 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5776 3488 5825 3516
rect 5776 3476 5782 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8444 3488 8953 3516
rect 8444 3476 8450 3488
rect 8941 3485 8953 3488
rect 8987 3516 8999 3519
rect 9582 3516 9588 3528
rect 8987 3488 9588 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 12710 3476 12716 3528
rect 12768 3476 12774 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13219 3488 13308 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 4448 3420 4554 3448
rect 3513 3383 3571 3389
rect 3513 3349 3525 3383
rect 3559 3380 3571 3383
rect 4448 3380 4476 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 6972 3420 7021 3448
rect 6972 3408 6978 3420
rect 7009 3417 7021 3420
rect 7055 3417 7067 3451
rect 7009 3411 7067 3417
rect 8018 3408 8024 3460
rect 8076 3408 8082 3460
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3417 8815 3451
rect 11606 3448 11612 3460
rect 11454 3420 11612 3448
rect 8757 3411 8815 3417
rect 3559 3352 4476 3380
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 6457 3383 6515 3389
rect 6457 3380 6469 3383
rect 6420 3352 6469 3380
rect 6420 3340 6426 3352
rect 6457 3349 6469 3352
rect 6503 3349 6515 3383
rect 6457 3343 6515 3349
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8772 3380 8800 3411
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 13280 3448 13308 3488
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 13556 3525 13584 3556
rect 15565 3553 15577 3556
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 16850 3584 16856 3596
rect 15979 3556 16856 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 16850 3544 16856 3556
rect 16908 3584 16914 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 16908 3556 18061 3584
rect 16908 3544 16914 3556
rect 18049 3553 18061 3556
rect 18095 3584 18107 3587
rect 19058 3584 19064 3596
rect 18095 3556 19064 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18380 3488 18613 3516
rect 18380 3476 18386 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 12584 3420 13308 3448
rect 12584 3408 12590 3420
rect 7432 3352 8800 3380
rect 7432 3340 7438 3352
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9180 3352 9229 3380
rect 9180 3340 9186 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 13280 3380 13308 3420
rect 13446 3408 13452 3460
rect 13504 3448 13510 3460
rect 14366 3448 14372 3460
rect 13504 3420 14372 3448
rect 13504 3408 13510 3420
rect 14366 3408 14372 3420
rect 14424 3408 14430 3460
rect 14826 3408 14832 3460
rect 14884 3408 14890 3460
rect 17342 3420 17448 3448
rect 14090 3380 14096 3392
rect 13280 3352 14096 3380
rect 9217 3343 9275 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 17420 3380 17448 3420
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17420 3352 18245 3380
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 18506 3340 18512 3392
rect 18564 3340 18570 3392
rect 1104 3290 26864 3312
rect 1104 3238 4829 3290
rect 4881 3238 4893 3290
rect 4945 3238 4957 3290
rect 5009 3238 5021 3290
rect 5073 3238 5085 3290
rect 5137 3238 11268 3290
rect 11320 3238 11332 3290
rect 11384 3238 11396 3290
rect 11448 3238 11460 3290
rect 11512 3238 11524 3290
rect 11576 3238 17707 3290
rect 17759 3238 17771 3290
rect 17823 3238 17835 3290
rect 17887 3238 17899 3290
rect 17951 3238 17963 3290
rect 18015 3238 24146 3290
rect 24198 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 26864 3290
rect 1104 3216 26864 3238
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6052 3148 6684 3176
rect 6052 3136 6058 3148
rect 4062 3108 4068 3120
rect 3712 3080 4068 3108
rect 3712 3049 3740 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4614 3068 4620 3120
rect 4672 3068 4678 3120
rect 6012 3049 6040 3136
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6236 3080 6561 3108
rect 6236 3068 6242 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6656 3108 6684 3148
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8018 3176 8024 3188
rect 7975 3148 8024 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8478 3136 8484 3188
rect 8536 3136 8542 3188
rect 8846 3136 8852 3188
rect 8904 3136 8910 3188
rect 10827 3179 10885 3185
rect 10827 3145 10839 3179
rect 10873 3176 10885 3179
rect 11054 3176 11060 3188
rect 10873 3148 11060 3176
rect 10873 3145 10885 3148
rect 10827 3139 10885 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 14826 3136 14832 3188
rect 14884 3136 14890 3188
rect 18414 3136 18420 3188
rect 18472 3136 18478 3188
rect 9122 3108 9128 3120
rect 6656 3080 7420 3108
rect 6549 3071 6607 3077
rect 7392 3052 7420 3080
rect 8588 3080 9128 3108
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 6779 3012 7052 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 3970 2932 3976 2984
rect 4028 2932 4034 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 5810 2972 5816 2984
rect 5675 2944 5816 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6270 2972 6276 2984
rect 6135 2944 6276 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7024 2981 7052 3012
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3040 8079 3043
rect 8386 3040 8392 3052
rect 8067 3012 8392 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 8588 3049 8616 3080
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 9766 3068 9772 3120
rect 9824 3068 9830 3120
rect 16850 3108 16856 3120
rect 16684 3080 16856 3108
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8720 3012 8769 3040
rect 8720 3000 8726 3012
rect 8757 3009 8769 3012
rect 8803 3040 8815 3043
rect 8938 3040 8944 3052
rect 8803 3012 8944 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3040 14979 3043
rect 15194 3040 15200 3052
rect 14967 3012 15200 3040
rect 14967 3009 14979 3012
rect 14921 3003 14979 3009
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 16684 3049 16712 3080
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 16942 3068 16948 3120
rect 17000 3068 17006 3120
rect 18506 3108 18512 3120
rect 18170 3080 18512 3108
rect 18506 3068 18512 3080
rect 18564 3068 18570 3120
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 7300 2904 7328 2935
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8352 2944 9045 2972
rect 8352 2932 8358 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 9950 2972 9956 2984
rect 9447 2944 9956 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 5592 2876 7328 2904
rect 5592 2864 5598 2876
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5718 2836 5724 2848
rect 5491 2808 5724 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5718 2796 5724 2808
rect 5776 2836 5782 2848
rect 6546 2836 6552 2848
rect 5776 2808 6552 2836
rect 5776 2796 5782 2808
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 1104 2746 26864 2768
rect 1104 2694 4169 2746
rect 4221 2694 4233 2746
rect 4285 2694 4297 2746
rect 4349 2694 4361 2746
rect 4413 2694 4425 2746
rect 4477 2694 10608 2746
rect 10660 2694 10672 2746
rect 10724 2694 10736 2746
rect 10788 2694 10800 2746
rect 10852 2694 10864 2746
rect 10916 2694 17047 2746
rect 17099 2694 17111 2746
rect 17163 2694 17175 2746
rect 17227 2694 17239 2746
rect 17291 2694 17303 2746
rect 17355 2694 23486 2746
rect 23538 2694 23550 2746
rect 23602 2694 23614 2746
rect 23666 2694 23678 2746
rect 23730 2694 23742 2746
rect 23794 2694 26864 2746
rect 1104 2672 26864 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2406 2632 2412 2644
rect 1627 2604 2412 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5592 2604 5733 2632
rect 5592 2592 5598 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 5721 2595 5779 2601
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 9766 2632 9772 2644
rect 9631 2604 9772 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10134 2496 10140 2508
rect 6748 2468 10140 2496
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6638 2428 6644 2440
rect 5951 2400 6644 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6748 2437 6776 2468
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 16356 2468 26004 2496
rect 16356 2456 16362 2468
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 8996 2400 9505 2428
rect 8996 2388 9002 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 11146 2428 11152 2440
rect 10459 2400 11152 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 14274 2388 14280 2440
rect 14332 2428 14338 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14332 2400 14473 2428
rect 14332 2388 14338 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 15838 2388 15844 2440
rect 15896 2428 15902 2440
rect 25976 2437 26004 2468
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 15896 2400 18061 2428
rect 15896 2388 15902 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 25961 2431 26019 2437
rect 25961 2397 25973 2431
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 6365 2363 6423 2369
rect 6365 2360 6377 2363
rect 6052 2332 6377 2360
rect 6052 2320 6058 2332
rect 6365 2329 6377 2332
rect 6411 2329 6423 2363
rect 6365 2323 6423 2329
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 10045 2363 10103 2369
rect 10045 2360 10057 2363
rect 10008 2332 10057 2360
rect 10008 2320 10014 2332
rect 10045 2329 10057 2332
rect 10091 2329 10103 2363
rect 10045 2323 10103 2329
rect 13906 2320 13912 2372
rect 13964 2360 13970 2372
rect 14093 2363 14151 2369
rect 14093 2360 14105 2363
rect 13964 2332 14105 2360
rect 13964 2320 13970 2332
rect 14093 2329 14105 2332
rect 14139 2329 14151 2363
rect 14093 2323 14151 2329
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 22005 2363 22063 2369
rect 22005 2360 22017 2363
rect 16448 2332 22017 2360
rect 16448 2320 16454 2332
rect 22005 2329 22017 2332
rect 22051 2329 22063 2363
rect 22005 2323 22063 2329
rect 18138 2252 18144 2304
rect 18196 2252 18202 2304
rect 21818 2252 21824 2304
rect 21876 2292 21882 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21876 2264 22109 2292
rect 21876 2252 21882 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22097 2255 22155 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 1104 2202 26864 2224
rect 1104 2150 4829 2202
rect 4881 2150 4893 2202
rect 4945 2150 4957 2202
rect 5009 2150 5021 2202
rect 5073 2150 5085 2202
rect 5137 2150 11268 2202
rect 11320 2150 11332 2202
rect 11384 2150 11396 2202
rect 11448 2150 11460 2202
rect 11512 2150 11524 2202
rect 11576 2150 17707 2202
rect 17759 2150 17771 2202
rect 17823 2150 17835 2202
rect 17887 2150 17899 2202
rect 17951 2150 17963 2202
rect 18015 2150 24146 2202
rect 24198 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 4169 27718 4221 27770
rect 4233 27718 4285 27770
rect 4297 27718 4349 27770
rect 4361 27718 4413 27770
rect 4425 27718 4477 27770
rect 10608 27718 10660 27770
rect 10672 27718 10724 27770
rect 10736 27718 10788 27770
rect 10800 27718 10852 27770
rect 10864 27718 10916 27770
rect 17047 27718 17099 27770
rect 17111 27718 17163 27770
rect 17175 27718 17227 27770
rect 17239 27718 17291 27770
rect 17303 27718 17355 27770
rect 23486 27718 23538 27770
rect 23550 27718 23602 27770
rect 23614 27718 23666 27770
rect 23678 27718 23730 27770
rect 23742 27718 23794 27770
rect 3424 27548 3476 27600
rect 10416 27548 10468 27600
rect 17408 27548 17460 27600
rect 24860 27591 24912 27600
rect 24860 27557 24869 27591
rect 24869 27557 24903 27591
rect 24903 27557 24912 27591
rect 24860 27548 24912 27557
rect 5356 27344 5408 27396
rect 7012 27344 7064 27396
rect 7104 27387 7156 27396
rect 7104 27353 7113 27387
rect 7113 27353 7147 27387
rect 7147 27353 7156 27387
rect 7104 27344 7156 27353
rect 10416 27344 10468 27396
rect 16580 27344 16632 27396
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 4344 27276 4396 27328
rect 4829 27174 4881 27226
rect 4893 27174 4945 27226
rect 4957 27174 5009 27226
rect 5021 27174 5073 27226
rect 5085 27174 5137 27226
rect 11268 27174 11320 27226
rect 11332 27174 11384 27226
rect 11396 27174 11448 27226
rect 11460 27174 11512 27226
rect 11524 27174 11576 27226
rect 17707 27174 17759 27226
rect 17771 27174 17823 27226
rect 17835 27174 17887 27226
rect 17899 27174 17951 27226
rect 17963 27174 18015 27226
rect 24146 27174 24198 27226
rect 24210 27174 24262 27226
rect 24274 27174 24326 27226
rect 24338 27174 24390 27226
rect 24402 27174 24454 27226
rect 4160 27072 4212 27124
rect 3332 26936 3384 26988
rect 4344 27004 4396 27056
rect 6368 26936 6420 26988
rect 5264 26868 5316 26920
rect 6736 26868 6788 26920
rect 6920 26979 6972 26988
rect 6920 26945 6929 26979
rect 6929 26945 6963 26979
rect 6963 26945 6972 26979
rect 6920 26936 6972 26945
rect 7196 26979 7248 26988
rect 7196 26945 7205 26979
rect 7205 26945 7239 26979
rect 7239 26945 7248 26979
rect 7196 26936 7248 26945
rect 5448 26800 5500 26852
rect 9128 26936 9180 26988
rect 14832 27072 14884 27124
rect 11980 26936 12032 26988
rect 18972 27004 19024 27056
rect 12256 26868 12308 26920
rect 17500 26868 17552 26920
rect 19708 26911 19760 26920
rect 19708 26877 19717 26911
rect 19717 26877 19751 26911
rect 19751 26877 19760 26911
rect 19708 26868 19760 26877
rect 19984 26911 20036 26920
rect 19984 26877 19993 26911
rect 19993 26877 20027 26911
rect 20027 26877 20036 26911
rect 19984 26868 20036 26877
rect 3608 26732 3660 26784
rect 7288 26732 7340 26784
rect 10324 26775 10376 26784
rect 10324 26741 10333 26775
rect 10333 26741 10367 26775
rect 10367 26741 10376 26775
rect 10324 26732 10376 26741
rect 12072 26732 12124 26784
rect 12716 26775 12768 26784
rect 12716 26741 12725 26775
rect 12725 26741 12759 26775
rect 12759 26741 12768 26775
rect 12716 26732 12768 26741
rect 13084 26775 13136 26784
rect 13084 26741 13093 26775
rect 13093 26741 13127 26775
rect 13127 26741 13136 26775
rect 13084 26732 13136 26741
rect 16212 26732 16264 26784
rect 16856 26732 16908 26784
rect 18144 26732 18196 26784
rect 4169 26630 4221 26682
rect 4233 26630 4285 26682
rect 4297 26630 4349 26682
rect 4361 26630 4413 26682
rect 4425 26630 4477 26682
rect 10608 26630 10660 26682
rect 10672 26630 10724 26682
rect 10736 26630 10788 26682
rect 10800 26630 10852 26682
rect 10864 26630 10916 26682
rect 17047 26630 17099 26682
rect 17111 26630 17163 26682
rect 17175 26630 17227 26682
rect 17239 26630 17291 26682
rect 17303 26630 17355 26682
rect 23486 26630 23538 26682
rect 23550 26630 23602 26682
rect 23614 26630 23666 26682
rect 23678 26630 23730 26682
rect 23742 26630 23794 26682
rect 3792 26528 3844 26580
rect 5448 26528 5500 26580
rect 7196 26528 7248 26580
rect 14372 26528 14424 26580
rect 18972 26571 19024 26580
rect 18972 26537 18981 26571
rect 18981 26537 19015 26571
rect 19015 26537 19024 26571
rect 18972 26528 19024 26537
rect 3884 26460 3936 26512
rect 3332 26367 3384 26376
rect 3332 26333 3341 26367
rect 3341 26333 3375 26367
rect 3375 26333 3384 26367
rect 3332 26324 3384 26333
rect 3608 26367 3660 26376
rect 3608 26333 3617 26367
rect 3617 26333 3651 26367
rect 3651 26333 3660 26367
rect 3608 26324 3660 26333
rect 3792 26367 3844 26376
rect 3792 26333 3801 26367
rect 3801 26333 3835 26367
rect 3835 26333 3844 26367
rect 3792 26324 3844 26333
rect 8116 26460 8168 26512
rect 15844 26503 15896 26512
rect 15844 26469 15853 26503
rect 15853 26469 15887 26503
rect 15887 26469 15896 26503
rect 15844 26460 15896 26469
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 5172 26256 5224 26308
rect 6644 26392 6696 26444
rect 13452 26392 13504 26444
rect 7196 26324 7248 26376
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 10876 26367 10928 26376
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 10876 26324 10928 26333
rect 10968 26324 11020 26376
rect 12900 26324 12952 26376
rect 3148 26188 3200 26240
rect 7380 26188 7432 26240
rect 10324 26256 10376 26308
rect 11612 26299 11664 26308
rect 11612 26265 11621 26299
rect 11621 26265 11655 26299
rect 11655 26265 11664 26299
rect 11612 26256 11664 26265
rect 12072 26256 12124 26308
rect 13176 26256 13228 26308
rect 15752 26392 15804 26444
rect 16672 26392 16724 26444
rect 19984 26392 20036 26444
rect 26148 26435 26200 26444
rect 26148 26401 26157 26435
rect 26157 26401 26191 26435
rect 26191 26401 26200 26435
rect 26148 26392 26200 26401
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 14464 26324 14516 26376
rect 14832 26367 14884 26376
rect 14832 26333 14841 26367
rect 14841 26333 14875 26367
rect 14875 26333 14884 26367
rect 14832 26324 14884 26333
rect 16028 26324 16080 26376
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 16212 26256 16264 26308
rect 16856 26256 16908 26308
rect 25504 26367 25556 26376
rect 25504 26333 25513 26367
rect 25513 26333 25547 26367
rect 25547 26333 25556 26367
rect 25504 26324 25556 26333
rect 19432 26256 19484 26308
rect 19616 26256 19668 26308
rect 21272 26299 21324 26308
rect 21272 26265 21281 26299
rect 21281 26265 21315 26299
rect 21315 26265 21324 26299
rect 21272 26256 21324 26265
rect 10784 26188 10836 26240
rect 12440 26188 12492 26240
rect 13544 26188 13596 26240
rect 13820 26188 13872 26240
rect 14740 26231 14792 26240
rect 14740 26197 14749 26231
rect 14749 26197 14783 26231
rect 14783 26197 14792 26231
rect 14740 26188 14792 26197
rect 15752 26188 15804 26240
rect 18052 26188 18104 26240
rect 19340 26188 19392 26240
rect 4829 26086 4881 26138
rect 4893 26086 4945 26138
rect 4957 26086 5009 26138
rect 5021 26086 5073 26138
rect 5085 26086 5137 26138
rect 11268 26086 11320 26138
rect 11332 26086 11384 26138
rect 11396 26086 11448 26138
rect 11460 26086 11512 26138
rect 11524 26086 11576 26138
rect 17707 26086 17759 26138
rect 17771 26086 17823 26138
rect 17835 26086 17887 26138
rect 17899 26086 17951 26138
rect 17963 26086 18015 26138
rect 24146 26086 24198 26138
rect 24210 26086 24262 26138
rect 24274 26086 24326 26138
rect 24338 26086 24390 26138
rect 24402 26086 24454 26138
rect 5172 25984 5224 26036
rect 7196 25984 7248 26036
rect 11612 25984 11664 26036
rect 11704 25984 11756 26036
rect 12256 25984 12308 26036
rect 6460 25916 6512 25968
rect 7104 25916 7156 25968
rect 7380 25916 7432 25968
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 6000 25848 6052 25900
rect 7564 25848 7616 25900
rect 9680 25916 9732 25968
rect 10968 25916 11020 25968
rect 11980 25959 12032 25968
rect 2964 25780 3016 25832
rect 3884 25780 3936 25832
rect 7012 25712 7064 25764
rect 7380 25780 7432 25832
rect 10784 25848 10836 25900
rect 11980 25925 11989 25959
rect 11989 25925 12023 25959
rect 12023 25925 12032 25959
rect 11980 25916 12032 25925
rect 12164 25916 12216 25968
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 11796 25848 11848 25857
rect 10232 25780 10284 25832
rect 10968 25823 11020 25832
rect 10968 25789 10977 25823
rect 10977 25789 11011 25823
rect 11011 25789 11020 25823
rect 10968 25780 11020 25789
rect 11704 25780 11756 25832
rect 12348 25891 12400 25900
rect 12348 25857 12357 25891
rect 12357 25857 12391 25891
rect 12391 25857 12400 25891
rect 12348 25848 12400 25857
rect 12440 25848 12492 25900
rect 13820 25984 13872 26036
rect 17500 25984 17552 26036
rect 19616 26027 19668 26036
rect 19616 25993 19625 26027
rect 19625 25993 19659 26027
rect 19659 25993 19668 26027
rect 19616 25984 19668 25993
rect 14740 25916 14792 25968
rect 15844 25916 15896 25968
rect 18052 25916 18104 25968
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 15936 25891 15988 25900
rect 15936 25857 15945 25891
rect 15945 25857 15979 25891
rect 15979 25857 15988 25891
rect 15936 25848 15988 25857
rect 16028 25891 16080 25900
rect 16028 25857 16037 25891
rect 16037 25857 16071 25891
rect 16071 25857 16080 25891
rect 16028 25848 16080 25857
rect 11980 25780 12032 25832
rect 12072 25780 12124 25832
rect 13360 25823 13412 25832
rect 13360 25789 13369 25823
rect 13369 25789 13403 25823
rect 13403 25789 13412 25823
rect 13360 25780 13412 25789
rect 13544 25780 13596 25832
rect 11520 25712 11572 25764
rect 12900 25712 12952 25764
rect 19340 25848 19392 25900
rect 20168 25848 20220 25900
rect 16672 25823 16724 25832
rect 16672 25789 16681 25823
rect 16681 25789 16715 25823
rect 16715 25789 16724 25823
rect 16672 25780 16724 25789
rect 5264 25644 5316 25696
rect 6920 25644 6972 25696
rect 11060 25644 11112 25696
rect 12992 25644 13044 25696
rect 14096 25644 14148 25696
rect 14556 25644 14608 25696
rect 17408 25644 17460 25696
rect 4169 25542 4221 25594
rect 4233 25542 4285 25594
rect 4297 25542 4349 25594
rect 4361 25542 4413 25594
rect 4425 25542 4477 25594
rect 10608 25542 10660 25594
rect 10672 25542 10724 25594
rect 10736 25542 10788 25594
rect 10800 25542 10852 25594
rect 10864 25542 10916 25594
rect 17047 25542 17099 25594
rect 17111 25542 17163 25594
rect 17175 25542 17227 25594
rect 17239 25542 17291 25594
rect 17303 25542 17355 25594
rect 23486 25542 23538 25594
rect 23550 25542 23602 25594
rect 23614 25542 23666 25594
rect 23678 25542 23730 25594
rect 23742 25542 23794 25594
rect 4528 25440 4580 25492
rect 7104 25483 7156 25492
rect 7104 25449 7113 25483
rect 7113 25449 7147 25483
rect 7147 25449 7156 25483
rect 7104 25440 7156 25449
rect 9680 25440 9732 25492
rect 11520 25483 11572 25492
rect 11520 25449 11529 25483
rect 11529 25449 11563 25483
rect 11563 25449 11572 25483
rect 11520 25440 11572 25449
rect 5448 25372 5500 25424
rect 6000 25372 6052 25424
rect 9128 25372 9180 25424
rect 12072 25440 12124 25492
rect 12164 25440 12216 25492
rect 13176 25440 13228 25492
rect 13360 25440 13412 25492
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 12348 25372 12400 25424
rect 13912 25483 13964 25492
rect 13912 25449 13921 25483
rect 13921 25449 13955 25483
rect 13955 25449 13964 25483
rect 13912 25440 13964 25449
rect 14464 25440 14516 25492
rect 16028 25440 16080 25492
rect 19708 25440 19760 25492
rect 16672 25372 16724 25424
rect 16948 25372 17000 25424
rect 18512 25372 18564 25424
rect 4528 25236 4580 25288
rect 5264 25236 5316 25288
rect 3608 25168 3660 25220
rect 4712 25168 4764 25220
rect 7656 25236 7708 25288
rect 13728 25304 13780 25356
rect 14372 25347 14424 25356
rect 14372 25313 14381 25347
rect 14381 25313 14415 25347
rect 14415 25313 14424 25347
rect 14372 25304 14424 25313
rect 10968 25236 11020 25288
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 4344 25143 4396 25152
rect 4344 25109 4353 25143
rect 4353 25109 4387 25143
rect 4387 25109 4396 25143
rect 4344 25100 4396 25109
rect 4620 25143 4672 25152
rect 4620 25109 4647 25143
rect 4647 25109 4672 25143
rect 4620 25100 4672 25109
rect 5172 25100 5224 25152
rect 6828 25100 6880 25152
rect 7196 25168 7248 25220
rect 7380 25168 7432 25220
rect 11888 25168 11940 25220
rect 10232 25143 10284 25152
rect 10232 25109 10241 25143
rect 10241 25109 10275 25143
rect 10275 25109 10284 25143
rect 10232 25100 10284 25109
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 13544 25236 13596 25288
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 14556 25279 14608 25288
rect 14556 25245 14565 25279
rect 14565 25245 14599 25279
rect 14599 25245 14608 25279
rect 14556 25236 14608 25245
rect 15200 25236 15252 25288
rect 15108 25211 15160 25220
rect 15108 25177 15117 25211
rect 15117 25177 15151 25211
rect 15151 25177 15160 25211
rect 15108 25168 15160 25177
rect 15660 25168 15712 25220
rect 16212 25279 16264 25288
rect 16212 25245 16221 25279
rect 16221 25245 16255 25279
rect 16255 25245 16264 25279
rect 16212 25236 16264 25245
rect 19340 25279 19392 25288
rect 19340 25245 19349 25279
rect 19349 25245 19383 25279
rect 19383 25245 19392 25279
rect 19340 25236 19392 25245
rect 16396 25211 16448 25220
rect 16396 25177 16405 25211
rect 16405 25177 16439 25211
rect 16439 25177 16448 25211
rect 16396 25168 16448 25177
rect 12440 25100 12492 25152
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 15752 25100 15804 25152
rect 18604 25168 18656 25220
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 19616 25279 19668 25288
rect 19616 25245 19625 25279
rect 19625 25245 19659 25279
rect 19659 25245 19668 25279
rect 19616 25236 19668 25245
rect 16856 25100 16908 25152
rect 18788 25100 18840 25152
rect 4829 24998 4881 25050
rect 4893 24998 4945 25050
rect 4957 24998 5009 25050
rect 5021 24998 5073 25050
rect 5085 24998 5137 25050
rect 11268 24998 11320 25050
rect 11332 24998 11384 25050
rect 11396 24998 11448 25050
rect 11460 24998 11512 25050
rect 11524 24998 11576 25050
rect 17707 24998 17759 25050
rect 17771 24998 17823 25050
rect 17835 24998 17887 25050
rect 17899 24998 17951 25050
rect 17963 24998 18015 25050
rect 24146 24998 24198 25050
rect 24210 24998 24262 25050
rect 24274 24998 24326 25050
rect 24338 24998 24390 25050
rect 24402 24998 24454 25050
rect 4436 24896 4488 24948
rect 6736 24896 6788 24948
rect 11796 24896 11848 24948
rect 11980 24896 12032 24948
rect 12808 24896 12860 24948
rect 13544 24896 13596 24948
rect 3148 24828 3200 24880
rect 4344 24828 4396 24880
rect 4620 24828 4672 24880
rect 5080 24828 5132 24880
rect 1400 24760 1452 24812
rect 3976 24803 4028 24812
rect 3976 24769 3985 24803
rect 3985 24769 4019 24803
rect 4019 24769 4028 24803
rect 3976 24760 4028 24769
rect 4068 24760 4120 24812
rect 2964 24692 3016 24744
rect 3884 24735 3936 24744
rect 3884 24701 3893 24735
rect 3893 24701 3927 24735
rect 3927 24701 3936 24735
rect 3884 24692 3936 24701
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 4804 24760 4856 24769
rect 5172 24760 5224 24812
rect 5264 24760 5316 24812
rect 5080 24692 5132 24744
rect 5540 24735 5592 24744
rect 5540 24701 5549 24735
rect 5549 24701 5583 24735
rect 5583 24701 5592 24735
rect 5540 24692 5592 24701
rect 5632 24735 5684 24744
rect 5632 24701 5641 24735
rect 5641 24701 5675 24735
rect 5675 24701 5684 24735
rect 5632 24692 5684 24701
rect 3608 24556 3660 24608
rect 3700 24599 3752 24608
rect 3700 24565 3709 24599
rect 3709 24565 3743 24599
rect 3743 24565 3752 24599
rect 3700 24556 3752 24565
rect 6184 24803 6236 24812
rect 6184 24769 6193 24803
rect 6193 24769 6227 24803
rect 6227 24769 6236 24803
rect 6184 24760 6236 24769
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 11704 24828 11756 24880
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 7012 24692 7064 24744
rect 8024 24735 8076 24744
rect 8024 24701 8033 24735
rect 8033 24701 8067 24735
rect 8067 24701 8076 24735
rect 8024 24692 8076 24701
rect 8116 24735 8168 24744
rect 8116 24701 8125 24735
rect 8125 24701 8159 24735
rect 8159 24701 8168 24735
rect 8116 24692 8168 24701
rect 8208 24735 8260 24744
rect 8208 24701 8217 24735
rect 8217 24701 8251 24735
rect 8251 24701 8260 24735
rect 8208 24692 8260 24701
rect 13820 24828 13872 24880
rect 14556 24896 14608 24948
rect 16396 24896 16448 24948
rect 14464 24828 14516 24880
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 12532 24692 12584 24744
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13452 24803 13504 24812
rect 13452 24769 13461 24803
rect 13461 24769 13495 24803
rect 13495 24769 13504 24803
rect 13452 24760 13504 24769
rect 15660 24828 15712 24880
rect 15936 24871 15988 24880
rect 15936 24837 15945 24871
rect 15945 24837 15979 24871
rect 15979 24837 15988 24871
rect 15936 24828 15988 24837
rect 14096 24692 14148 24744
rect 15108 24692 15160 24744
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18604 24760 18656 24812
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 18972 24803 19024 24812
rect 18972 24769 18989 24803
rect 18989 24769 19024 24803
rect 18972 24760 19024 24769
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 19432 24803 19484 24812
rect 19432 24769 19441 24803
rect 19441 24769 19475 24803
rect 19475 24769 19484 24803
rect 19432 24760 19484 24769
rect 19616 24828 19668 24880
rect 19892 24828 19944 24880
rect 6736 24556 6788 24608
rect 7104 24556 7156 24608
rect 12256 24624 12308 24676
rect 13176 24624 13228 24676
rect 7748 24599 7800 24608
rect 7748 24565 7757 24599
rect 7757 24565 7791 24599
rect 7791 24565 7800 24599
rect 7748 24556 7800 24565
rect 12440 24556 12492 24608
rect 13084 24556 13136 24608
rect 13912 24556 13964 24608
rect 19340 24624 19392 24676
rect 19800 24735 19852 24744
rect 19800 24701 19809 24735
rect 19809 24701 19843 24735
rect 19843 24701 19852 24735
rect 19800 24692 19852 24701
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 21272 24828 21324 24880
rect 22560 24828 22612 24880
rect 20076 24760 20128 24769
rect 21640 24692 21692 24744
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 18512 24556 18564 24608
rect 19156 24556 19208 24608
rect 23296 24556 23348 24608
rect 4169 24454 4221 24506
rect 4233 24454 4285 24506
rect 4297 24454 4349 24506
rect 4361 24454 4413 24506
rect 4425 24454 4477 24506
rect 10608 24454 10660 24506
rect 10672 24454 10724 24506
rect 10736 24454 10788 24506
rect 10800 24454 10852 24506
rect 10864 24454 10916 24506
rect 17047 24454 17099 24506
rect 17111 24454 17163 24506
rect 17175 24454 17227 24506
rect 17239 24454 17291 24506
rect 17303 24454 17355 24506
rect 23486 24454 23538 24506
rect 23550 24454 23602 24506
rect 23614 24454 23666 24506
rect 23678 24454 23730 24506
rect 23742 24454 23794 24506
rect 3148 24352 3200 24404
rect 3884 24352 3936 24404
rect 4068 24327 4120 24336
rect 4068 24293 4077 24327
rect 4077 24293 4111 24327
rect 4111 24293 4120 24327
rect 4068 24284 4120 24293
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 3700 24216 3752 24268
rect 4528 24216 4580 24268
rect 4804 24352 4856 24404
rect 5540 24352 5592 24404
rect 6552 24352 6604 24404
rect 7012 24352 7064 24404
rect 7656 24352 7708 24404
rect 12900 24352 12952 24404
rect 13268 24352 13320 24404
rect 15936 24352 15988 24404
rect 18972 24352 19024 24404
rect 19432 24352 19484 24404
rect 22560 24352 22612 24404
rect 6184 24284 6236 24336
rect 11060 24284 11112 24336
rect 18604 24284 18656 24336
rect 19340 24284 19392 24336
rect 20076 24284 20128 24336
rect 22192 24284 22244 24336
rect 2872 24148 2924 24200
rect 3608 24148 3660 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4252 24191 4304 24200
rect 4252 24157 4261 24191
rect 4261 24157 4295 24191
rect 4295 24157 4304 24191
rect 4252 24148 4304 24157
rect 2780 24080 2832 24132
rect 4620 24080 4672 24132
rect 4804 24148 4856 24200
rect 5448 24148 5500 24200
rect 7748 24216 7800 24268
rect 18512 24216 18564 24268
rect 7104 24148 7156 24200
rect 7380 24148 7432 24200
rect 8208 24148 8260 24200
rect 13728 24148 13780 24200
rect 19156 24148 19208 24200
rect 20444 24216 20496 24268
rect 23296 24259 23348 24268
rect 23296 24225 23305 24259
rect 23305 24225 23339 24259
rect 23339 24225 23348 24259
rect 23296 24216 23348 24225
rect 10692 24080 10744 24132
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 12992 24080 13044 24089
rect 13176 24123 13228 24132
rect 13176 24089 13201 24123
rect 13201 24089 13228 24123
rect 13176 24080 13228 24089
rect 19248 24080 19300 24132
rect 21272 24148 21324 24200
rect 20628 24080 20680 24132
rect 22652 24148 22704 24200
rect 4252 24012 4304 24064
rect 5632 24012 5684 24064
rect 6828 24012 6880 24064
rect 9956 24012 10008 24064
rect 13544 24055 13596 24064
rect 13544 24021 13553 24055
rect 13553 24021 13587 24055
rect 13587 24021 13596 24055
rect 13544 24012 13596 24021
rect 21916 24012 21968 24064
rect 4829 23910 4881 23962
rect 4893 23910 4945 23962
rect 4957 23910 5009 23962
rect 5021 23910 5073 23962
rect 5085 23910 5137 23962
rect 11268 23910 11320 23962
rect 11332 23910 11384 23962
rect 11396 23910 11448 23962
rect 11460 23910 11512 23962
rect 11524 23910 11576 23962
rect 17707 23910 17759 23962
rect 17771 23910 17823 23962
rect 17835 23910 17887 23962
rect 17899 23910 17951 23962
rect 17963 23910 18015 23962
rect 24146 23910 24198 23962
rect 24210 23910 24262 23962
rect 24274 23910 24326 23962
rect 24338 23910 24390 23962
rect 24402 23910 24454 23962
rect 2780 23851 2832 23860
rect 2780 23817 2789 23851
rect 2789 23817 2823 23851
rect 2823 23817 2832 23851
rect 2780 23808 2832 23817
rect 3976 23808 4028 23860
rect 5540 23808 5592 23860
rect 940 23672 992 23724
rect 2872 23715 2924 23724
rect 2872 23681 2881 23715
rect 2881 23681 2915 23715
rect 2915 23681 2924 23715
rect 2872 23672 2924 23681
rect 4252 23740 4304 23792
rect 7104 23740 7156 23792
rect 8208 23808 8260 23860
rect 9312 23740 9364 23792
rect 4620 23672 4672 23724
rect 6276 23672 6328 23724
rect 6644 23672 6696 23724
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 10232 23808 10284 23860
rect 10508 23808 10560 23860
rect 13820 23808 13872 23860
rect 19800 23851 19852 23860
rect 19800 23817 19809 23851
rect 19809 23817 19843 23851
rect 19843 23817 19852 23851
rect 19800 23808 19852 23817
rect 13084 23740 13136 23792
rect 10324 23715 10376 23724
rect 10324 23681 10342 23715
rect 10342 23681 10376 23715
rect 10324 23672 10376 23681
rect 4160 23647 4212 23656
rect 4160 23613 4169 23647
rect 4169 23613 4203 23647
rect 4203 23613 4212 23647
rect 4160 23604 4212 23613
rect 4712 23604 4764 23656
rect 9772 23604 9824 23656
rect 9956 23604 10008 23656
rect 11704 23672 11756 23724
rect 12624 23672 12676 23724
rect 13544 23672 13596 23724
rect 13820 23672 13872 23724
rect 18236 23740 18288 23792
rect 19156 23740 19208 23792
rect 14832 23672 14884 23724
rect 10600 23604 10652 23656
rect 5264 23536 5316 23588
rect 2780 23468 2832 23520
rect 9680 23468 9732 23520
rect 10692 23579 10744 23588
rect 10692 23545 10701 23579
rect 10701 23545 10735 23579
rect 10735 23545 10744 23579
rect 15200 23647 15252 23656
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 10692 23536 10744 23545
rect 10968 23468 11020 23520
rect 12072 23468 12124 23520
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14372 23468 14424 23520
rect 16304 23511 16356 23520
rect 16304 23477 16313 23511
rect 16313 23477 16347 23511
rect 16347 23477 16356 23511
rect 16304 23468 16356 23477
rect 19340 23672 19392 23724
rect 19892 23672 19944 23724
rect 20904 23672 20956 23724
rect 21916 23740 21968 23792
rect 22192 23808 22244 23860
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 21548 23672 21600 23724
rect 19340 23536 19392 23588
rect 20628 23604 20680 23656
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 22100 23468 22152 23520
rect 22284 23511 22336 23520
rect 22284 23477 22293 23511
rect 22293 23477 22327 23511
rect 22327 23477 22336 23511
rect 22284 23468 22336 23477
rect 22652 23468 22704 23520
rect 4169 23366 4221 23418
rect 4233 23366 4285 23418
rect 4297 23366 4349 23418
rect 4361 23366 4413 23418
rect 4425 23366 4477 23418
rect 10608 23366 10660 23418
rect 10672 23366 10724 23418
rect 10736 23366 10788 23418
rect 10800 23366 10852 23418
rect 10864 23366 10916 23418
rect 17047 23366 17099 23418
rect 17111 23366 17163 23418
rect 17175 23366 17227 23418
rect 17239 23366 17291 23418
rect 17303 23366 17355 23418
rect 23486 23366 23538 23418
rect 23550 23366 23602 23418
rect 23614 23366 23666 23418
rect 23678 23366 23730 23418
rect 23742 23366 23794 23418
rect 7104 23307 7156 23316
rect 7104 23273 7113 23307
rect 7113 23273 7147 23307
rect 7147 23273 7156 23307
rect 7104 23264 7156 23273
rect 9128 23264 9180 23316
rect 9404 23264 9456 23316
rect 8116 23196 8168 23248
rect 8944 23196 8996 23248
rect 2872 23128 2924 23180
rect 2780 23103 2832 23112
rect 2780 23069 2789 23103
rect 2789 23069 2823 23103
rect 2823 23069 2832 23103
rect 2780 23060 2832 23069
rect 3240 23060 3292 23112
rect 6184 23060 6236 23112
rect 6736 23128 6788 23180
rect 9036 23128 9088 23180
rect 9588 23171 9640 23180
rect 9588 23137 9597 23171
rect 9597 23137 9631 23171
rect 9631 23137 9640 23171
rect 9588 23128 9640 23137
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 10508 23264 10560 23316
rect 7104 23060 7156 23112
rect 8392 23060 8444 23112
rect 9772 23103 9824 23112
rect 9772 23069 9790 23103
rect 9790 23069 9824 23103
rect 9772 23060 9824 23069
rect 10508 23128 10560 23180
rect 12440 23264 12492 23316
rect 12808 23264 12860 23316
rect 15660 23264 15712 23316
rect 19708 23264 19760 23316
rect 19892 23307 19944 23316
rect 19892 23273 19901 23307
rect 19901 23273 19935 23307
rect 19935 23273 19944 23307
rect 19892 23264 19944 23273
rect 20076 23307 20128 23316
rect 20076 23273 20085 23307
rect 20085 23273 20119 23307
rect 20119 23273 20128 23307
rect 20076 23264 20128 23273
rect 20904 23307 20956 23316
rect 20904 23273 20913 23307
rect 20913 23273 20947 23307
rect 20947 23273 20956 23307
rect 20904 23264 20956 23273
rect 11796 23196 11848 23248
rect 12992 23196 13044 23248
rect 12164 23128 12216 23180
rect 10692 23060 10744 23112
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 11428 23103 11480 23112
rect 11428 23069 11437 23103
rect 11437 23069 11471 23103
rect 11471 23069 11480 23103
rect 11428 23060 11480 23069
rect 11704 23060 11756 23112
rect 11888 23060 11940 23112
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 14188 23128 14240 23180
rect 16672 23128 16724 23180
rect 6000 23035 6052 23044
rect 6000 23001 6009 23035
rect 6009 23001 6043 23035
rect 6043 23001 6052 23035
rect 6000 22992 6052 23001
rect 8024 22992 8076 23044
rect 13820 23060 13872 23112
rect 16856 23103 16908 23112
rect 16856 23069 16865 23103
rect 16865 23069 16899 23103
rect 16899 23069 16908 23103
rect 16856 23060 16908 23069
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 19340 23196 19392 23248
rect 19064 23103 19116 23112
rect 19064 23069 19073 23103
rect 19073 23069 19107 23103
rect 19107 23069 19116 23103
rect 19064 23060 19116 23069
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 19708 23060 19760 23112
rect 8852 22924 8904 22976
rect 10232 22924 10284 22976
rect 11612 22924 11664 22976
rect 12072 22924 12124 22976
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 12900 22967 12952 22976
rect 12900 22933 12909 22967
rect 12909 22933 12943 22967
rect 12943 22933 12952 22967
rect 12900 22924 12952 22933
rect 13268 22992 13320 23044
rect 16304 22992 16356 23044
rect 20444 23060 20496 23112
rect 19892 22992 19944 23044
rect 20536 23035 20588 23044
rect 13452 22924 13504 22976
rect 19616 22924 19668 22976
rect 19800 22967 19852 22976
rect 19800 22933 19809 22967
rect 19809 22933 19843 22967
rect 19843 22933 19852 22967
rect 19800 22924 19852 22933
rect 20536 23001 20563 23035
rect 20563 23001 20588 23035
rect 20536 22992 20588 23001
rect 20720 23035 20772 23044
rect 20720 23001 20729 23035
rect 20729 23001 20763 23035
rect 20763 23001 20772 23035
rect 20720 22992 20772 23001
rect 22100 23264 22152 23316
rect 22284 23128 22336 23180
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 21272 23035 21324 23044
rect 21272 23001 21281 23035
rect 21281 23001 21315 23035
rect 21315 23001 21324 23035
rect 21272 22992 21324 23001
rect 20812 22924 20864 22976
rect 22100 22924 22152 22976
rect 22652 22992 22704 23044
rect 4829 22822 4881 22874
rect 4893 22822 4945 22874
rect 4957 22822 5009 22874
rect 5021 22822 5073 22874
rect 5085 22822 5137 22874
rect 11268 22822 11320 22874
rect 11332 22822 11384 22874
rect 11396 22822 11448 22874
rect 11460 22822 11512 22874
rect 11524 22822 11576 22874
rect 17707 22822 17759 22874
rect 17771 22822 17823 22874
rect 17835 22822 17887 22874
rect 17899 22822 17951 22874
rect 17963 22822 18015 22874
rect 24146 22822 24198 22874
rect 24210 22822 24262 22874
rect 24274 22822 24326 22874
rect 24338 22822 24390 22874
rect 24402 22822 24454 22874
rect 6552 22720 6604 22772
rect 8208 22652 8260 22704
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 8852 22584 8904 22636
rect 11520 22720 11572 22772
rect 11888 22720 11940 22772
rect 11980 22720 12032 22772
rect 9680 22627 9732 22636
rect 9680 22593 9689 22627
rect 9689 22593 9723 22627
rect 9723 22593 9732 22627
rect 9680 22584 9732 22593
rect 9220 22559 9272 22568
rect 9220 22525 9229 22559
rect 9229 22525 9263 22559
rect 9263 22525 9272 22559
rect 9220 22516 9272 22525
rect 9496 22516 9548 22568
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 9128 22380 9180 22432
rect 9864 22448 9916 22500
rect 10140 22584 10192 22636
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 11060 22559 11112 22568
rect 11060 22525 11069 22559
rect 11069 22525 11103 22559
rect 11103 22525 11112 22559
rect 11060 22516 11112 22525
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 12440 22652 12492 22704
rect 13452 22720 13504 22772
rect 15200 22720 15252 22772
rect 16948 22720 17000 22772
rect 12256 22516 12308 22568
rect 12440 22516 12492 22568
rect 12900 22584 12952 22636
rect 14372 22652 14424 22704
rect 17960 22652 18012 22704
rect 19984 22652 20036 22704
rect 13360 22584 13412 22636
rect 13820 22627 13872 22636
rect 13820 22593 13829 22627
rect 13829 22593 13863 22627
rect 13863 22593 13872 22627
rect 13820 22584 13872 22593
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 21640 22652 21692 22704
rect 20628 22627 20680 22636
rect 20628 22593 20637 22627
rect 20637 22593 20671 22627
rect 20671 22593 20680 22627
rect 20628 22584 20680 22593
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 22100 22695 22152 22704
rect 22100 22661 22109 22695
rect 22109 22661 22143 22695
rect 22143 22661 22152 22695
rect 22100 22652 22152 22661
rect 22652 22652 22704 22704
rect 14188 22516 14240 22568
rect 16580 22516 16632 22568
rect 12992 22448 13044 22500
rect 18604 22516 18656 22568
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 19708 22516 19760 22568
rect 19800 22516 19852 22568
rect 20536 22448 20588 22500
rect 21548 22516 21600 22568
rect 21640 22516 21692 22568
rect 10048 22380 10100 22432
rect 10416 22380 10468 22432
rect 10692 22380 10744 22432
rect 11336 22380 11388 22432
rect 11888 22380 11940 22432
rect 12256 22380 12308 22432
rect 13268 22423 13320 22432
rect 13268 22389 13277 22423
rect 13277 22389 13311 22423
rect 13311 22389 13320 22423
rect 13268 22380 13320 22389
rect 14648 22380 14700 22432
rect 16764 22380 16816 22432
rect 20720 22380 20772 22432
rect 21548 22380 21600 22432
rect 4169 22278 4221 22330
rect 4233 22278 4285 22330
rect 4297 22278 4349 22330
rect 4361 22278 4413 22330
rect 4425 22278 4477 22330
rect 10608 22278 10660 22330
rect 10672 22278 10724 22330
rect 10736 22278 10788 22330
rect 10800 22278 10852 22330
rect 10864 22278 10916 22330
rect 17047 22278 17099 22330
rect 17111 22278 17163 22330
rect 17175 22278 17227 22330
rect 17239 22278 17291 22330
rect 17303 22278 17355 22330
rect 23486 22278 23538 22330
rect 23550 22278 23602 22330
rect 23614 22278 23666 22330
rect 23678 22278 23730 22330
rect 23742 22278 23794 22330
rect 4344 22176 4396 22228
rect 4712 22176 4764 22228
rect 9128 22219 9180 22228
rect 9128 22185 9137 22219
rect 9137 22185 9171 22219
rect 9171 22185 9180 22219
rect 9128 22176 9180 22185
rect 9864 22176 9916 22228
rect 9956 22219 10008 22228
rect 9956 22185 9965 22219
rect 9965 22185 9999 22219
rect 9999 22185 10008 22219
rect 9956 22176 10008 22185
rect 10324 22176 10376 22228
rect 10600 22176 10652 22228
rect 11152 22176 11204 22228
rect 11336 22176 11388 22228
rect 12440 22176 12492 22228
rect 12532 22176 12584 22228
rect 13268 22176 13320 22228
rect 14188 22219 14240 22228
rect 14188 22185 14197 22219
rect 14197 22185 14231 22219
rect 14231 22185 14240 22219
rect 14188 22176 14240 22185
rect 16580 22176 16632 22228
rect 16764 22176 16816 22228
rect 18512 22219 18564 22228
rect 18512 22185 18521 22219
rect 18521 22185 18555 22219
rect 18555 22185 18564 22219
rect 18512 22176 18564 22185
rect 18972 22219 19024 22228
rect 18972 22185 18981 22219
rect 18981 22185 19015 22219
rect 19015 22185 19024 22219
rect 18972 22176 19024 22185
rect 19064 22176 19116 22228
rect 940 21972 992 22024
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 2872 22015 2924 22024
rect 2412 21972 2464 21981
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 2504 21879 2556 21888
rect 2504 21845 2513 21879
rect 2513 21845 2547 21879
rect 2547 21845 2556 21879
rect 2504 21836 2556 21845
rect 2780 21879 2832 21888
rect 2780 21845 2789 21879
rect 2789 21845 2823 21879
rect 2823 21845 2832 21879
rect 2780 21836 2832 21845
rect 2964 21879 3016 21888
rect 2964 21845 2973 21879
rect 2973 21845 3007 21879
rect 3007 21845 3016 21879
rect 2964 21836 3016 21845
rect 3332 22015 3384 22024
rect 3332 21981 3341 22015
rect 3341 21981 3375 22015
rect 3375 21981 3384 22015
rect 3332 21972 3384 21981
rect 9496 22108 9548 22160
rect 11612 22108 11664 22160
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 4160 22015 4212 22024
rect 4160 21981 4169 22015
rect 4169 21981 4203 22015
rect 4203 21981 4212 22015
rect 4160 21972 4212 21981
rect 3516 21904 3568 21956
rect 3700 21836 3752 21888
rect 5080 21972 5132 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 6276 22040 6328 22092
rect 9128 22040 9180 22092
rect 5448 21904 5500 21956
rect 4436 21879 4488 21888
rect 4436 21845 4445 21879
rect 4445 21845 4479 21879
rect 4479 21845 4488 21879
rect 4436 21836 4488 21845
rect 4712 21836 4764 21888
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 5356 21836 5408 21888
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 8392 21972 8444 22024
rect 9404 22015 9456 22024
rect 6184 21947 6236 21956
rect 6184 21913 6193 21947
rect 6193 21913 6227 21947
rect 6227 21913 6236 21947
rect 6184 21904 6236 21913
rect 7196 21904 7248 21956
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 9956 21972 10008 22024
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 12072 22108 12124 22160
rect 20076 22176 20128 22228
rect 20536 22219 20588 22228
rect 20536 22185 20545 22219
rect 20545 22185 20579 22219
rect 20579 22185 20588 22219
rect 20536 22176 20588 22185
rect 21364 22176 21416 22228
rect 11612 21972 11664 21981
rect 9496 21904 9548 21956
rect 9864 21904 9916 21956
rect 6460 21836 6512 21888
rect 6828 21836 6880 21888
rect 9680 21836 9732 21888
rect 10232 21904 10284 21956
rect 10508 21904 10560 21956
rect 16396 22040 16448 22092
rect 16856 22040 16908 22092
rect 17960 22040 18012 22092
rect 21640 22108 21692 22160
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 10140 21879 10192 21888
rect 10140 21845 10149 21879
rect 10149 21845 10183 21879
rect 10183 21845 10192 21879
rect 10140 21836 10192 21845
rect 10968 21836 11020 21888
rect 15200 21904 15252 21956
rect 15660 21947 15712 21956
rect 15660 21913 15669 21947
rect 15669 21913 15703 21947
rect 15703 21913 15712 21947
rect 15660 21904 15712 21913
rect 16764 21972 16816 22024
rect 17592 21972 17644 22024
rect 18052 21972 18104 22024
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 19892 22040 19944 22092
rect 20812 22040 20864 22092
rect 21548 22083 21600 22092
rect 21548 22049 21557 22083
rect 21557 22049 21591 22083
rect 21591 22049 21600 22083
rect 21548 22040 21600 22049
rect 22652 22083 22704 22092
rect 22652 22049 22661 22083
rect 22661 22049 22695 22083
rect 22695 22049 22704 22083
rect 22652 22040 22704 22049
rect 18604 21904 18656 21956
rect 20076 22015 20128 22024
rect 20076 21981 20085 22015
rect 20085 21981 20119 22015
rect 20119 21981 20128 22015
rect 20076 21972 20128 21981
rect 20628 21972 20680 22024
rect 21640 22015 21692 22024
rect 21640 21981 21649 22015
rect 21649 21981 21683 22015
rect 21683 21981 21692 22015
rect 21640 21972 21692 21981
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 18236 21836 18288 21888
rect 18696 21836 18748 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 20076 21836 20128 21888
rect 4829 21734 4881 21786
rect 4893 21734 4945 21786
rect 4957 21734 5009 21786
rect 5021 21734 5073 21786
rect 5085 21734 5137 21786
rect 11268 21734 11320 21786
rect 11332 21734 11384 21786
rect 11396 21734 11448 21786
rect 11460 21734 11512 21786
rect 11524 21734 11576 21786
rect 17707 21734 17759 21786
rect 17771 21734 17823 21786
rect 17835 21734 17887 21786
rect 17899 21734 17951 21786
rect 17963 21734 18015 21786
rect 24146 21734 24198 21786
rect 24210 21734 24262 21786
rect 24274 21734 24326 21786
rect 24338 21734 24390 21786
rect 24402 21734 24454 21786
rect 3332 21632 3384 21684
rect 3792 21632 3844 21684
rect 3516 21564 3568 21616
rect 6184 21632 6236 21684
rect 6460 21675 6512 21684
rect 6460 21641 6469 21675
rect 6469 21641 6503 21675
rect 6503 21641 6512 21675
rect 6460 21632 6512 21641
rect 7196 21632 7248 21684
rect 8208 21632 8260 21684
rect 10232 21632 10284 21684
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 15200 21632 15252 21684
rect 15660 21675 15712 21684
rect 15660 21641 15669 21675
rect 15669 21641 15703 21675
rect 15703 21641 15712 21675
rect 15660 21632 15712 21641
rect 18328 21632 18380 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2780 21496 2832 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4712 21564 4764 21616
rect 3884 21428 3936 21480
rect 4344 21428 4396 21480
rect 4712 21428 4764 21480
rect 5172 21505 5181 21538
rect 5181 21505 5215 21538
rect 5215 21505 5224 21538
rect 5172 21486 5224 21505
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 12440 21564 12492 21616
rect 13544 21564 13596 21616
rect 5724 21496 5776 21548
rect 6828 21496 6880 21548
rect 7104 21496 7156 21548
rect 15936 21564 15988 21616
rect 16764 21564 16816 21616
rect 14464 21496 14516 21548
rect 15292 21496 15344 21548
rect 6000 21471 6052 21480
rect 6000 21437 6009 21471
rect 6009 21437 6043 21471
rect 6043 21437 6052 21471
rect 6000 21428 6052 21437
rect 6552 21428 6604 21480
rect 6460 21360 6512 21412
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 16396 21496 16448 21548
rect 18972 21564 19024 21616
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 17592 21428 17644 21480
rect 20076 21428 20128 21480
rect 3792 21292 3844 21344
rect 4344 21292 4396 21344
rect 4896 21292 4948 21344
rect 5356 21292 5408 21344
rect 5632 21335 5684 21344
rect 5632 21301 5641 21335
rect 5641 21301 5675 21335
rect 5675 21301 5684 21335
rect 5632 21292 5684 21301
rect 5816 21292 5868 21344
rect 6828 21335 6880 21344
rect 6828 21301 6837 21335
rect 6837 21301 6871 21335
rect 6871 21301 6880 21335
rect 6828 21292 6880 21301
rect 13268 21292 13320 21344
rect 18788 21292 18840 21344
rect 4169 21190 4221 21242
rect 4233 21190 4285 21242
rect 4297 21190 4349 21242
rect 4361 21190 4413 21242
rect 4425 21190 4477 21242
rect 10608 21190 10660 21242
rect 10672 21190 10724 21242
rect 10736 21190 10788 21242
rect 10800 21190 10852 21242
rect 10864 21190 10916 21242
rect 17047 21190 17099 21242
rect 17111 21190 17163 21242
rect 17175 21190 17227 21242
rect 17239 21190 17291 21242
rect 17303 21190 17355 21242
rect 23486 21190 23538 21242
rect 23550 21190 23602 21242
rect 23614 21190 23666 21242
rect 23678 21190 23730 21242
rect 23742 21190 23794 21242
rect 3884 21131 3936 21140
rect 3884 21097 3893 21131
rect 3893 21097 3927 21131
rect 3927 21097 3936 21131
rect 3884 21088 3936 21097
rect 4896 21088 4948 21140
rect 5172 21131 5224 21140
rect 5172 21097 5181 21131
rect 5181 21097 5215 21131
rect 5215 21097 5224 21131
rect 5172 21088 5224 21097
rect 5356 21088 5408 21140
rect 9956 21088 10008 21140
rect 14004 21088 14056 21140
rect 16948 21131 17000 21140
rect 16948 21097 16957 21131
rect 16957 21097 16991 21131
rect 16991 21097 17000 21131
rect 16948 21088 17000 21097
rect 1400 20952 1452 21004
rect 2964 20952 3016 21004
rect 4160 21020 4212 21072
rect 5264 21020 5316 21072
rect 10324 21020 10376 21072
rect 13544 21020 13596 21072
rect 5632 20952 5684 21004
rect 8944 20995 8996 21004
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 9404 20952 9456 21004
rect 2504 20816 2556 20868
rect 3792 20816 3844 20868
rect 4804 20927 4856 20936
rect 4804 20893 4813 20927
rect 4813 20893 4847 20927
rect 4847 20893 4856 20927
rect 4804 20884 4856 20893
rect 4620 20816 4672 20868
rect 5356 20884 5408 20936
rect 7012 20859 7064 20868
rect 7012 20825 7021 20859
rect 7021 20825 7055 20859
rect 7055 20825 7064 20859
rect 7012 20816 7064 20825
rect 9036 20816 9088 20868
rect 9680 20884 9732 20936
rect 13452 20952 13504 21004
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 10324 20884 10376 20936
rect 9956 20859 10008 20868
rect 9956 20825 9965 20859
rect 9965 20825 9999 20859
rect 9999 20825 10008 20859
rect 9956 20816 10008 20825
rect 15292 20884 15344 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 5908 20748 5960 20800
rect 6460 20748 6512 20800
rect 8668 20748 8720 20800
rect 9772 20791 9824 20800
rect 9772 20757 9781 20791
rect 9781 20757 9815 20791
rect 9815 20757 9824 20791
rect 9772 20748 9824 20757
rect 9864 20748 9916 20800
rect 14464 20859 14516 20868
rect 14464 20825 14473 20859
rect 14473 20825 14507 20859
rect 14507 20825 14516 20859
rect 14464 20816 14516 20825
rect 15108 20816 15160 20868
rect 15660 20859 15712 20868
rect 15660 20825 15669 20859
rect 15669 20825 15703 20859
rect 15703 20825 15712 20859
rect 15660 20816 15712 20825
rect 17408 20748 17460 20800
rect 4829 20646 4881 20698
rect 4893 20646 4945 20698
rect 4957 20646 5009 20698
rect 5021 20646 5073 20698
rect 5085 20646 5137 20698
rect 11268 20646 11320 20698
rect 11332 20646 11384 20698
rect 11396 20646 11448 20698
rect 11460 20646 11512 20698
rect 11524 20646 11576 20698
rect 17707 20646 17759 20698
rect 17771 20646 17823 20698
rect 17835 20646 17887 20698
rect 17899 20646 17951 20698
rect 17963 20646 18015 20698
rect 24146 20646 24198 20698
rect 24210 20646 24262 20698
rect 24274 20646 24326 20698
rect 24338 20646 24390 20698
rect 24402 20646 24454 20698
rect 3516 20544 3568 20596
rect 3976 20544 4028 20596
rect 4712 20544 4764 20596
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 8208 20587 8260 20596
rect 3792 20476 3844 20528
rect 5172 20519 5224 20528
rect 5172 20485 5199 20519
rect 5199 20485 5224 20519
rect 5172 20476 5224 20485
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 5632 20476 5684 20528
rect 3700 20408 3752 20417
rect 4160 20340 4212 20392
rect 3608 20272 3660 20324
rect 4068 20272 4120 20324
rect 5724 20408 5776 20460
rect 6000 20408 6052 20460
rect 8208 20553 8217 20587
rect 8217 20553 8251 20587
rect 8251 20553 8260 20587
rect 8208 20544 8260 20553
rect 8944 20544 8996 20596
rect 9772 20544 9824 20596
rect 10048 20544 10100 20596
rect 7288 20476 7340 20528
rect 6460 20451 6512 20460
rect 6460 20417 6469 20451
rect 6469 20417 6503 20451
rect 6503 20417 6512 20451
rect 6460 20408 6512 20417
rect 9680 20408 9732 20460
rect 9956 20451 10008 20460
rect 5448 20272 5500 20324
rect 6736 20383 6788 20392
rect 6736 20349 6745 20383
rect 6745 20349 6779 20383
rect 6779 20349 6788 20383
rect 6736 20340 6788 20349
rect 9956 20417 9973 20451
rect 9973 20417 10008 20451
rect 9956 20408 10008 20417
rect 11336 20476 11388 20528
rect 11704 20544 11756 20596
rect 17040 20544 17092 20596
rect 24584 20544 24636 20596
rect 10876 20408 10928 20460
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 11796 20408 11848 20460
rect 17408 20476 17460 20528
rect 18604 20476 18656 20528
rect 18788 20476 18840 20528
rect 10508 20340 10560 20392
rect 10232 20272 10284 20324
rect 15384 20383 15436 20392
rect 15384 20349 15393 20383
rect 15393 20349 15427 20383
rect 15427 20349 15436 20383
rect 15384 20340 15436 20349
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16856 20408 16908 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 16488 20340 16540 20392
rect 14464 20272 14516 20324
rect 16396 20315 16448 20324
rect 16396 20281 16405 20315
rect 16405 20281 16439 20315
rect 16439 20281 16448 20315
rect 16396 20272 16448 20281
rect 16948 20272 17000 20324
rect 17500 20340 17552 20392
rect 17684 20340 17736 20392
rect 18420 20340 18472 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 4528 20204 4580 20256
rect 5632 20204 5684 20256
rect 5816 20204 5868 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 10324 20204 10376 20256
rect 11152 20204 11204 20256
rect 16120 20204 16172 20256
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 4169 20102 4221 20154
rect 4233 20102 4285 20154
rect 4297 20102 4349 20154
rect 4361 20102 4413 20154
rect 4425 20102 4477 20154
rect 10608 20102 10660 20154
rect 10672 20102 10724 20154
rect 10736 20102 10788 20154
rect 10800 20102 10852 20154
rect 10864 20102 10916 20154
rect 17047 20102 17099 20154
rect 17111 20102 17163 20154
rect 17175 20102 17227 20154
rect 17239 20102 17291 20154
rect 17303 20102 17355 20154
rect 23486 20102 23538 20154
rect 23550 20102 23602 20154
rect 23614 20102 23666 20154
rect 23678 20102 23730 20154
rect 23742 20102 23794 20154
rect 6736 20000 6788 20052
rect 7288 20043 7340 20052
rect 7288 20009 7297 20043
rect 7297 20009 7331 20043
rect 7331 20009 7340 20043
rect 7288 20000 7340 20009
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 9588 20000 9640 20052
rect 940 19796 992 19848
rect 4620 19796 4672 19848
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 5448 19796 5500 19848
rect 5540 19839 5592 19848
rect 5540 19805 5549 19839
rect 5549 19805 5583 19839
rect 5583 19805 5592 19839
rect 5540 19796 5592 19805
rect 5816 19796 5868 19848
rect 8392 19864 8444 19916
rect 7104 19796 7156 19848
rect 4712 19728 4764 19780
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 9864 19932 9916 19984
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 11152 19864 11204 19916
rect 8944 19728 8996 19780
rect 9496 19728 9548 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 3516 19660 3568 19712
rect 8760 19660 8812 19712
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10416 19796 10468 19848
rect 10876 19796 10928 19848
rect 11336 19839 11388 19848
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 11612 19864 11664 19916
rect 11612 19728 11664 19780
rect 16120 20043 16172 20052
rect 16120 20009 16129 20043
rect 16129 20009 16163 20043
rect 16163 20009 16172 20043
rect 16120 20000 16172 20009
rect 16488 20043 16540 20052
rect 16488 20009 16497 20043
rect 16497 20009 16531 20043
rect 16531 20009 16540 20043
rect 16488 20000 16540 20009
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 14464 19907 14516 19916
rect 14464 19873 14473 19907
rect 14473 19873 14507 19907
rect 14507 19873 14516 19907
rect 14464 19864 14516 19873
rect 16672 19864 16724 19916
rect 12808 19728 12860 19780
rect 11060 19660 11112 19712
rect 13728 19660 13780 19712
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 15844 19796 15896 19848
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 16396 19796 16448 19848
rect 17684 20000 17736 20052
rect 17500 19864 17552 19916
rect 18420 20043 18472 20052
rect 18420 20009 18429 20043
rect 18429 20009 18463 20043
rect 18463 20009 18472 20043
rect 18420 20000 18472 20009
rect 18604 20000 18656 20052
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 14924 19771 14976 19780
rect 14924 19737 14933 19771
rect 14933 19737 14967 19771
rect 14967 19737 14976 19771
rect 14924 19728 14976 19737
rect 17592 19796 17644 19848
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 19524 19864 19576 19916
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 18972 19796 19024 19848
rect 19156 19796 19208 19848
rect 18328 19728 18380 19780
rect 16028 19660 16080 19712
rect 18052 19660 18104 19712
rect 19984 19728 20036 19780
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 4829 19558 4881 19610
rect 4893 19558 4945 19610
rect 4957 19558 5009 19610
rect 5021 19558 5073 19610
rect 5085 19558 5137 19610
rect 11268 19558 11320 19610
rect 11332 19558 11384 19610
rect 11396 19558 11448 19610
rect 11460 19558 11512 19610
rect 11524 19558 11576 19610
rect 17707 19558 17759 19610
rect 17771 19558 17823 19610
rect 17835 19558 17887 19610
rect 17899 19558 17951 19610
rect 17963 19558 18015 19610
rect 24146 19558 24198 19610
rect 24210 19558 24262 19610
rect 24274 19558 24326 19610
rect 24338 19558 24390 19610
rect 24402 19558 24454 19610
rect 2872 19456 2924 19508
rect 4160 19456 4212 19508
rect 5356 19456 5408 19508
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 3332 19320 3384 19372
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 3884 19388 3936 19440
rect 4160 19320 4212 19372
rect 4528 19320 4580 19372
rect 3148 19252 3200 19304
rect 4804 19252 4856 19304
rect 3332 19184 3384 19236
rect 4068 19184 4120 19236
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 5724 19363 5776 19372
rect 5724 19329 5733 19363
rect 5733 19329 5767 19363
rect 5767 19329 5776 19363
rect 5724 19320 5776 19329
rect 9404 19456 9456 19508
rect 10416 19456 10468 19508
rect 10600 19456 10652 19508
rect 6920 19388 6972 19440
rect 11612 19456 11664 19508
rect 16488 19456 16540 19508
rect 6276 19320 6328 19372
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9220 19320 9272 19372
rect 13728 19431 13780 19440
rect 13728 19397 13737 19431
rect 13737 19397 13771 19431
rect 13771 19397 13780 19431
rect 13728 19388 13780 19397
rect 16580 19388 16632 19440
rect 16948 19456 17000 19508
rect 16764 19388 16816 19440
rect 19156 19456 19208 19508
rect 19524 19456 19576 19508
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 9588 19320 9640 19372
rect 10048 19320 10100 19372
rect 10600 19320 10652 19372
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 11152 19320 11204 19372
rect 11796 19320 11848 19372
rect 12532 19320 12584 19372
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 6736 19252 6788 19304
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 10232 19184 10284 19236
rect 10876 19252 10928 19304
rect 11704 19252 11756 19304
rect 16488 19363 16540 19372
rect 16488 19329 16497 19363
rect 16497 19329 16531 19363
rect 16531 19329 16540 19363
rect 16488 19320 16540 19329
rect 18880 19388 18932 19440
rect 20444 19388 20496 19440
rect 11060 19184 11112 19236
rect 11888 19184 11940 19236
rect 15476 19184 15528 19236
rect 15936 19184 15988 19236
rect 16764 19252 16816 19304
rect 16396 19184 16448 19236
rect 18052 19252 18104 19304
rect 20076 19252 20128 19304
rect 12808 19116 12860 19168
rect 14188 19116 14240 19168
rect 16764 19116 16816 19168
rect 16856 19116 16908 19168
rect 18604 19116 18656 19168
rect 4169 19014 4221 19066
rect 4233 19014 4285 19066
rect 4297 19014 4349 19066
rect 4361 19014 4413 19066
rect 4425 19014 4477 19066
rect 10608 19014 10660 19066
rect 10672 19014 10724 19066
rect 10736 19014 10788 19066
rect 10800 19014 10852 19066
rect 10864 19014 10916 19066
rect 17047 19014 17099 19066
rect 17111 19014 17163 19066
rect 17175 19014 17227 19066
rect 17239 19014 17291 19066
rect 17303 19014 17355 19066
rect 23486 19014 23538 19066
rect 23550 19014 23602 19066
rect 23614 19014 23666 19066
rect 23678 19014 23730 19066
rect 23742 19014 23794 19066
rect 5724 18912 5776 18964
rect 6920 18955 6972 18964
rect 6920 18921 6929 18955
rect 6929 18921 6963 18955
rect 6963 18921 6972 18955
rect 6920 18912 6972 18921
rect 9036 18912 9088 18964
rect 10232 18912 10284 18964
rect 10508 18912 10560 18964
rect 12532 18955 12584 18964
rect 12532 18921 12541 18955
rect 12541 18921 12575 18955
rect 12575 18921 12584 18955
rect 12532 18912 12584 18921
rect 15384 18912 15436 18964
rect 16212 18912 16264 18964
rect 17316 18912 17368 18964
rect 3148 18776 3200 18828
rect 3332 18776 3384 18828
rect 1492 18751 1544 18760
rect 1492 18717 1501 18751
rect 1501 18717 1535 18751
rect 1535 18717 1544 18751
rect 1492 18708 1544 18717
rect 2872 18708 2924 18760
rect 4620 18819 4672 18828
rect 4620 18785 4629 18819
rect 4629 18785 4663 18819
rect 4663 18785 4672 18819
rect 4620 18776 4672 18785
rect 4804 18776 4856 18828
rect 4528 18708 4580 18760
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 5448 18708 5500 18760
rect 7104 18844 7156 18896
rect 10416 18844 10468 18896
rect 8760 18708 8812 18760
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 9404 18708 9456 18760
rect 9588 18708 9640 18760
rect 11060 18776 11112 18828
rect 15936 18844 15988 18896
rect 16488 18844 16540 18896
rect 16764 18844 16816 18896
rect 14924 18776 14976 18828
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10508 18751 10560 18760
rect 10508 18717 10517 18751
rect 10517 18717 10551 18751
rect 10551 18717 10560 18751
rect 10508 18708 10560 18717
rect 5540 18640 5592 18692
rect 12808 18708 12860 18760
rect 3884 18615 3936 18624
rect 3884 18581 3893 18615
rect 3893 18581 3927 18615
rect 3927 18581 3936 18615
rect 3884 18572 3936 18581
rect 8300 18572 8352 18624
rect 10048 18572 10100 18624
rect 15108 18751 15160 18760
rect 15108 18717 15117 18751
rect 15117 18717 15151 18751
rect 15151 18717 15160 18751
rect 15108 18708 15160 18717
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 15476 18708 15528 18760
rect 15752 18708 15804 18760
rect 15568 18572 15620 18624
rect 15936 18683 15988 18692
rect 15936 18649 15945 18683
rect 15945 18649 15979 18683
rect 15979 18649 15988 18683
rect 15936 18640 15988 18649
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 16856 18708 16908 18760
rect 18144 18912 18196 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 20076 18955 20128 18964
rect 20076 18921 20085 18955
rect 20085 18921 20119 18955
rect 20119 18921 20128 18955
rect 20076 18912 20128 18921
rect 20444 18955 20496 18964
rect 20444 18921 20453 18955
rect 20453 18921 20487 18955
rect 20487 18921 20496 18955
rect 20444 18912 20496 18921
rect 18052 18776 18104 18828
rect 19800 18776 19852 18828
rect 17960 18708 18012 18760
rect 18604 18708 18656 18760
rect 18788 18708 18840 18760
rect 17408 18640 17460 18692
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 26516 18751 26568 18760
rect 26516 18717 26525 18751
rect 26525 18717 26559 18751
rect 26559 18717 26568 18751
rect 26516 18708 26568 18717
rect 16028 18572 16080 18624
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 17040 18572 17092 18624
rect 17684 18572 17736 18624
rect 18328 18572 18380 18624
rect 19432 18572 19484 18624
rect 4829 18470 4881 18522
rect 4893 18470 4945 18522
rect 4957 18470 5009 18522
rect 5021 18470 5073 18522
rect 5085 18470 5137 18522
rect 11268 18470 11320 18522
rect 11332 18470 11384 18522
rect 11396 18470 11448 18522
rect 11460 18470 11512 18522
rect 11524 18470 11576 18522
rect 17707 18470 17759 18522
rect 17771 18470 17823 18522
rect 17835 18470 17887 18522
rect 17899 18470 17951 18522
rect 17963 18470 18015 18522
rect 24146 18470 24198 18522
rect 24210 18470 24262 18522
rect 24274 18470 24326 18522
rect 24338 18470 24390 18522
rect 24402 18470 24454 18522
rect 2780 18368 2832 18420
rect 5172 18368 5224 18420
rect 10232 18368 10284 18420
rect 14556 18368 14608 18420
rect 15108 18368 15160 18420
rect 3884 18300 3936 18352
rect 1492 18232 1544 18284
rect 10232 18232 10284 18284
rect 10324 18232 10376 18284
rect 13728 18232 13780 18284
rect 12532 18164 12584 18216
rect 12716 18096 12768 18148
rect 13544 18164 13596 18216
rect 14188 18164 14240 18216
rect 14832 18207 14884 18216
rect 14832 18173 14841 18207
rect 14841 18173 14875 18207
rect 14875 18173 14884 18207
rect 14832 18164 14884 18173
rect 15568 18368 15620 18420
rect 16212 18368 16264 18420
rect 16948 18368 17000 18420
rect 17316 18368 17368 18420
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 15936 18232 15988 18284
rect 16856 18232 16908 18284
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 20996 18368 21048 18420
rect 19432 18343 19484 18352
rect 19432 18309 19441 18343
rect 19441 18309 19475 18343
rect 19475 18309 19484 18343
rect 19432 18300 19484 18309
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 16580 18096 16632 18148
rect 19340 18096 19392 18148
rect 15476 18028 15528 18080
rect 15936 18028 15988 18080
rect 16396 18028 16448 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 16948 18028 17000 18080
rect 18328 18028 18380 18080
rect 4169 17926 4221 17978
rect 4233 17926 4285 17978
rect 4297 17926 4349 17978
rect 4361 17926 4413 17978
rect 4425 17926 4477 17978
rect 10608 17926 10660 17978
rect 10672 17926 10724 17978
rect 10736 17926 10788 17978
rect 10800 17926 10852 17978
rect 10864 17926 10916 17978
rect 17047 17926 17099 17978
rect 17111 17926 17163 17978
rect 17175 17926 17227 17978
rect 17239 17926 17291 17978
rect 17303 17926 17355 17978
rect 23486 17926 23538 17978
rect 23550 17926 23602 17978
rect 23614 17926 23666 17978
rect 23678 17926 23730 17978
rect 23742 17926 23794 17978
rect 3424 17824 3476 17876
rect 6644 17824 6696 17876
rect 10048 17824 10100 17876
rect 11060 17824 11112 17876
rect 12716 17867 12768 17876
rect 12716 17833 12725 17867
rect 12725 17833 12759 17867
rect 12759 17833 12768 17867
rect 12716 17824 12768 17833
rect 13544 17824 13596 17876
rect 15476 17867 15528 17876
rect 15476 17833 15485 17867
rect 15485 17833 15519 17867
rect 15519 17833 15528 17867
rect 15476 17824 15528 17833
rect 16672 17824 16724 17876
rect 10692 17799 10744 17808
rect 10692 17765 10701 17799
rect 10701 17765 10735 17799
rect 10735 17765 10744 17799
rect 10692 17756 10744 17765
rect 10876 17756 10928 17808
rect 15752 17756 15804 17808
rect 940 17620 992 17672
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 9404 17620 9456 17672
rect 10324 17620 10376 17672
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 10692 17552 10744 17604
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 6276 17484 6328 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 10600 17527 10652 17536
rect 10600 17493 10609 17527
rect 10609 17493 10643 17527
rect 10643 17493 10652 17527
rect 10600 17484 10652 17493
rect 11152 17484 11204 17536
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14004 17620 14056 17672
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 18144 17620 18196 17672
rect 21824 17620 21876 17672
rect 19064 17484 19116 17536
rect 21640 17552 21692 17604
rect 4829 17382 4881 17434
rect 4893 17382 4945 17434
rect 4957 17382 5009 17434
rect 5021 17382 5073 17434
rect 5085 17382 5137 17434
rect 11268 17382 11320 17434
rect 11332 17382 11384 17434
rect 11396 17382 11448 17434
rect 11460 17382 11512 17434
rect 11524 17382 11576 17434
rect 17707 17382 17759 17434
rect 17771 17382 17823 17434
rect 17835 17382 17887 17434
rect 17899 17382 17951 17434
rect 17963 17382 18015 17434
rect 24146 17382 24198 17434
rect 24210 17382 24262 17434
rect 24274 17382 24326 17434
rect 24338 17382 24390 17434
rect 24402 17382 24454 17434
rect 1584 17280 1636 17332
rect 3884 17144 3936 17196
rect 4068 16940 4120 16992
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 5080 17187 5132 17196
rect 5080 17153 5114 17187
rect 5114 17153 5132 17187
rect 5080 17144 5132 17153
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11152 17280 11204 17332
rect 9772 17255 9824 17264
rect 9772 17221 9781 17255
rect 9781 17221 9815 17255
rect 9815 17221 9824 17255
rect 9772 17212 9824 17221
rect 8300 17144 8352 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 10600 17144 10652 17196
rect 14096 17212 14148 17264
rect 14832 17280 14884 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 19340 17280 19392 17332
rect 13728 17144 13780 17196
rect 6276 17076 6328 17128
rect 8484 17119 8536 17128
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 8576 17008 8628 17060
rect 9220 17076 9272 17128
rect 10508 17076 10560 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11612 17076 11664 17128
rect 15292 17212 15344 17264
rect 17960 17212 18012 17264
rect 16764 17144 16816 17196
rect 18236 17144 18288 17196
rect 19156 17212 19208 17264
rect 10140 17008 10192 17060
rect 11244 17008 11296 17060
rect 5540 16940 5592 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 11060 16940 11112 16992
rect 11796 16940 11848 16992
rect 15660 17119 15712 17128
rect 15660 17085 15669 17119
rect 15669 17085 15703 17119
rect 15703 17085 15712 17119
rect 15660 17076 15712 17085
rect 12808 16940 12860 16992
rect 13636 17008 13688 17060
rect 15844 17008 15896 17060
rect 18328 17008 18380 17060
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 22928 17144 22980 17196
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 19064 17119 19116 17128
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 18788 17008 18840 17060
rect 13728 16940 13780 16992
rect 14004 16940 14056 16992
rect 15752 16983 15804 16992
rect 15752 16949 15761 16983
rect 15761 16949 15795 16983
rect 15795 16949 15804 16983
rect 15752 16940 15804 16949
rect 16672 16940 16724 16992
rect 18236 16940 18288 16992
rect 19248 16940 19300 16992
rect 22100 16940 22152 16992
rect 4169 16838 4221 16890
rect 4233 16838 4285 16890
rect 4297 16838 4349 16890
rect 4361 16838 4413 16890
rect 4425 16838 4477 16890
rect 10608 16838 10660 16890
rect 10672 16838 10724 16890
rect 10736 16838 10788 16890
rect 10800 16838 10852 16890
rect 10864 16838 10916 16890
rect 17047 16838 17099 16890
rect 17111 16838 17163 16890
rect 17175 16838 17227 16890
rect 17239 16838 17291 16890
rect 17303 16838 17355 16890
rect 23486 16838 23538 16890
rect 23550 16838 23602 16890
rect 23614 16838 23666 16890
rect 23678 16838 23730 16890
rect 23742 16838 23794 16890
rect 1492 16600 1544 16652
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 4804 16736 4856 16788
rect 5080 16736 5132 16788
rect 5540 16736 5592 16788
rect 8300 16736 8352 16788
rect 8484 16736 8536 16788
rect 9220 16736 9272 16788
rect 4068 16575 4120 16584
rect 4068 16541 4102 16575
rect 4102 16541 4120 16575
rect 4068 16532 4120 16541
rect 5080 16532 5132 16584
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 8576 16668 8628 16720
rect 9404 16668 9456 16720
rect 9864 16736 9916 16788
rect 8484 16600 8536 16652
rect 9772 16600 9824 16652
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 11244 16736 11296 16788
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 13544 16736 13596 16788
rect 15752 16736 15804 16788
rect 17040 16779 17092 16788
rect 17040 16745 17049 16779
rect 17049 16745 17083 16779
rect 17083 16745 17092 16779
rect 17040 16736 17092 16745
rect 17960 16736 18012 16788
rect 18420 16736 18472 16788
rect 18696 16736 18748 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 11612 16600 11664 16652
rect 15200 16668 15252 16720
rect 12348 16575 12400 16584
rect 2228 16464 2280 16516
rect 2872 16396 2924 16448
rect 3792 16464 3844 16516
rect 6552 16507 6604 16516
rect 6552 16473 6586 16507
rect 6586 16473 6604 16507
rect 6552 16464 6604 16473
rect 6644 16464 6696 16516
rect 11060 16464 11112 16516
rect 11336 16464 11388 16516
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 12348 16532 12400 16541
rect 12900 16532 12952 16584
rect 14740 16532 14792 16584
rect 18972 16668 19024 16720
rect 19248 16668 19300 16720
rect 16580 16600 16632 16652
rect 18420 16600 18472 16652
rect 18788 16600 18840 16652
rect 16764 16532 16816 16584
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 5080 16396 5132 16448
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 7288 16396 7340 16448
rect 7748 16396 7800 16448
rect 10968 16396 11020 16448
rect 11704 16396 11756 16448
rect 11888 16439 11940 16448
rect 11888 16405 11897 16439
rect 11897 16405 11931 16439
rect 11931 16405 11940 16439
rect 11888 16396 11940 16405
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 12348 16396 12400 16448
rect 14280 16396 14332 16448
rect 14832 16396 14884 16448
rect 16856 16464 16908 16516
rect 16948 16464 17000 16516
rect 18236 16532 18288 16584
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 18512 16532 18564 16584
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 21364 16532 21416 16584
rect 22928 16736 22980 16788
rect 23020 16736 23072 16788
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 17592 16396 17644 16448
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 21640 16464 21692 16516
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 23848 16668 23900 16720
rect 22284 16464 22336 16516
rect 18328 16396 18380 16448
rect 19800 16439 19852 16448
rect 19800 16405 19809 16439
rect 19809 16405 19843 16439
rect 19843 16405 19852 16439
rect 19800 16396 19852 16405
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 22468 16439 22520 16448
rect 22468 16405 22477 16439
rect 22477 16405 22511 16439
rect 22511 16405 22520 16439
rect 22468 16396 22520 16405
rect 23204 16396 23256 16448
rect 24032 16575 24084 16584
rect 24032 16541 24041 16575
rect 24041 16541 24075 16575
rect 24075 16541 24084 16575
rect 24032 16532 24084 16541
rect 24032 16396 24084 16448
rect 4829 16294 4881 16346
rect 4893 16294 4945 16346
rect 4957 16294 5009 16346
rect 5021 16294 5073 16346
rect 5085 16294 5137 16346
rect 11268 16294 11320 16346
rect 11332 16294 11384 16346
rect 11396 16294 11448 16346
rect 11460 16294 11512 16346
rect 11524 16294 11576 16346
rect 17707 16294 17759 16346
rect 17771 16294 17823 16346
rect 17835 16294 17887 16346
rect 17899 16294 17951 16346
rect 17963 16294 18015 16346
rect 24146 16294 24198 16346
rect 24210 16294 24262 16346
rect 24274 16294 24326 16346
rect 24338 16294 24390 16346
rect 24402 16294 24454 16346
rect 6552 16192 6604 16244
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 8392 16192 8444 16244
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 9956 16235 10008 16244
rect 9956 16201 9965 16235
rect 9965 16201 9999 16235
rect 9999 16201 10008 16235
rect 9956 16192 10008 16201
rect 3976 16124 4028 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 5172 16056 5224 16108
rect 5724 16056 5776 16108
rect 6276 16124 6328 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7196 16124 7248 16176
rect 7288 16167 7340 16176
rect 7288 16133 7297 16167
rect 7297 16133 7331 16167
rect 7331 16133 7340 16167
rect 7288 16124 7340 16133
rect 7380 16124 7432 16176
rect 8576 16056 8628 16108
rect 11888 16192 11940 16244
rect 14096 16192 14148 16244
rect 14280 16235 14332 16244
rect 14280 16201 14289 16235
rect 14289 16201 14323 16235
rect 14323 16201 14332 16235
rect 14280 16192 14332 16201
rect 14648 16192 14700 16244
rect 7748 15988 7800 16040
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 11612 16056 11664 16108
rect 12348 16124 12400 16176
rect 13084 16124 13136 16176
rect 17960 16192 18012 16244
rect 16672 16124 16724 16176
rect 16948 16124 17000 16176
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 17592 16124 17644 16176
rect 16580 16056 16632 16108
rect 18328 16124 18380 16176
rect 23940 16235 23992 16244
rect 23940 16201 23949 16235
rect 23949 16201 23983 16235
rect 23983 16201 23992 16235
rect 23940 16192 23992 16201
rect 20352 16124 20404 16176
rect 21364 16124 21416 16176
rect 4068 15920 4120 15972
rect 6920 15920 6972 15972
rect 7288 15920 7340 15972
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 12348 16031 12400 16040
rect 12348 15997 12357 16031
rect 12357 15997 12391 16031
rect 12391 15997 12400 16031
rect 12348 15988 12400 15997
rect 3424 15852 3476 15904
rect 3608 15852 3660 15904
rect 4528 15852 4580 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 7380 15852 7432 15904
rect 7656 15852 7708 15904
rect 7748 15852 7800 15904
rect 10140 15895 10192 15904
rect 10140 15861 10149 15895
rect 10149 15861 10183 15895
rect 10183 15861 10192 15895
rect 10140 15852 10192 15861
rect 10508 15852 10560 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 16764 15988 16816 16040
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18420 16056 18472 16108
rect 18972 16056 19024 16108
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 21824 16099 21876 16108
rect 21824 16065 21833 16099
rect 21833 16065 21867 16099
rect 21867 16065 21876 16099
rect 21824 16056 21876 16065
rect 22468 16124 22520 16176
rect 17408 15920 17460 15972
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 16948 15852 17000 15904
rect 18144 15988 18196 16040
rect 19340 16031 19392 16040
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 20720 15988 20772 16040
rect 22836 15988 22888 16040
rect 24032 16099 24084 16108
rect 24032 16065 24041 16099
rect 24041 16065 24075 16099
rect 24075 16065 24084 16099
rect 24032 16056 24084 16065
rect 24584 16056 24636 16108
rect 25044 16056 25096 16108
rect 24492 15920 24544 15972
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 22560 15852 22612 15904
rect 23204 15895 23256 15904
rect 23204 15861 23213 15895
rect 23213 15861 23247 15895
rect 23247 15861 23256 15895
rect 23204 15852 23256 15861
rect 23388 15852 23440 15904
rect 25136 15895 25188 15904
rect 25136 15861 25145 15895
rect 25145 15861 25179 15895
rect 25179 15861 25188 15895
rect 25136 15852 25188 15861
rect 4169 15750 4221 15802
rect 4233 15750 4285 15802
rect 4297 15750 4349 15802
rect 4361 15750 4413 15802
rect 4425 15750 4477 15802
rect 10608 15750 10660 15802
rect 10672 15750 10724 15802
rect 10736 15750 10788 15802
rect 10800 15750 10852 15802
rect 10864 15750 10916 15802
rect 17047 15750 17099 15802
rect 17111 15750 17163 15802
rect 17175 15750 17227 15802
rect 17239 15750 17291 15802
rect 17303 15750 17355 15802
rect 23486 15750 23538 15802
rect 23550 15750 23602 15802
rect 23614 15750 23666 15802
rect 23678 15750 23730 15802
rect 23742 15750 23794 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2228 15648 2280 15700
rect 3148 15648 3200 15700
rect 3608 15691 3660 15700
rect 3608 15657 3617 15691
rect 3617 15657 3651 15691
rect 3651 15657 3660 15691
rect 3608 15648 3660 15657
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 8484 15648 8536 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 11612 15648 11664 15700
rect 12348 15648 12400 15700
rect 13084 15691 13136 15700
rect 13084 15657 13093 15691
rect 13093 15657 13127 15691
rect 13127 15657 13136 15691
rect 13084 15648 13136 15657
rect 15016 15691 15068 15700
rect 15016 15657 15025 15691
rect 15025 15657 15059 15691
rect 15059 15657 15068 15691
rect 15016 15648 15068 15657
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 17500 15691 17552 15700
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17500 15648 17552 15657
rect 19340 15648 19392 15700
rect 21640 15691 21692 15700
rect 21640 15657 21649 15691
rect 21649 15657 21683 15691
rect 21683 15657 21692 15691
rect 21640 15648 21692 15657
rect 21824 15648 21876 15700
rect 2872 15580 2924 15632
rect 4620 15580 4672 15632
rect 3332 15512 3384 15564
rect 3884 15512 3936 15564
rect 4068 15512 4120 15564
rect 4344 15512 4396 15564
rect 16856 15580 16908 15632
rect 18052 15580 18104 15632
rect 18328 15580 18380 15632
rect 22284 15580 22336 15632
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 3424 15444 3476 15453
rect 4528 15444 4580 15496
rect 6552 15512 6604 15564
rect 6276 15444 6328 15496
rect 2780 15351 2832 15360
rect 2780 15317 2789 15351
rect 2789 15317 2823 15351
rect 2823 15317 2832 15351
rect 2780 15308 2832 15317
rect 5632 15376 5684 15428
rect 7288 15444 7340 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 9680 15512 9732 15564
rect 10048 15512 10100 15564
rect 12072 15512 12124 15564
rect 8484 15444 8536 15496
rect 13912 15512 13964 15564
rect 13176 15444 13228 15496
rect 14740 15444 14792 15496
rect 16948 15512 17000 15564
rect 17960 15512 18012 15564
rect 18788 15512 18840 15564
rect 20996 15512 21048 15564
rect 15476 15444 15528 15496
rect 16304 15444 16356 15496
rect 18420 15444 18472 15496
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 3332 15308 3384 15360
rect 10508 15419 10560 15428
rect 10508 15385 10517 15419
rect 10517 15385 10551 15419
rect 10551 15385 10560 15419
rect 10508 15376 10560 15385
rect 11244 15376 11296 15428
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 7380 15308 7432 15360
rect 7748 15308 7800 15360
rect 16488 15376 16540 15428
rect 16672 15376 16724 15428
rect 18052 15376 18104 15428
rect 19064 15376 19116 15428
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 22100 15444 22152 15496
rect 23388 15444 23440 15496
rect 24032 15487 24084 15496
rect 24032 15453 24041 15487
rect 24041 15453 24075 15487
rect 24075 15453 24084 15487
rect 24032 15444 24084 15453
rect 25136 15444 25188 15496
rect 18328 15308 18380 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 20996 15376 21048 15428
rect 21364 15419 21416 15428
rect 21364 15385 21373 15419
rect 21373 15385 21407 15419
rect 21407 15385 21416 15419
rect 21364 15376 21416 15385
rect 19800 15308 19852 15317
rect 20904 15351 20956 15360
rect 20904 15317 20913 15351
rect 20913 15317 20947 15351
rect 20947 15317 20956 15351
rect 20904 15308 20956 15317
rect 22836 15308 22888 15360
rect 22928 15308 22980 15360
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 4829 15206 4881 15258
rect 4893 15206 4945 15258
rect 4957 15206 5009 15258
rect 5021 15206 5073 15258
rect 5085 15206 5137 15258
rect 11268 15206 11320 15258
rect 11332 15206 11384 15258
rect 11396 15206 11448 15258
rect 11460 15206 11512 15258
rect 11524 15206 11576 15258
rect 17707 15206 17759 15258
rect 17771 15206 17823 15258
rect 17835 15206 17887 15258
rect 17899 15206 17951 15258
rect 17963 15206 18015 15258
rect 24146 15206 24198 15258
rect 24210 15206 24262 15258
rect 24274 15206 24326 15258
rect 24338 15206 24390 15258
rect 24402 15206 24454 15258
rect 2780 15104 2832 15156
rect 3148 15104 3200 15156
rect 3976 15104 4028 15156
rect 5724 15104 5776 15156
rect 3056 15079 3108 15088
rect 3056 15045 3065 15079
rect 3065 15045 3099 15079
rect 3099 15045 3108 15079
rect 3056 15036 3108 15045
rect 3792 15036 3844 15088
rect 4068 15036 4120 15088
rect 16580 15104 16632 15156
rect 16672 15147 16724 15156
rect 16672 15113 16681 15147
rect 16681 15113 16715 15147
rect 16715 15113 16724 15147
rect 16672 15104 16724 15113
rect 18236 15104 18288 15156
rect 6644 14968 6696 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 16764 15036 16816 15088
rect 16948 15036 17000 15088
rect 6920 14900 6972 14952
rect 7288 14900 7340 14952
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 18144 14968 18196 15020
rect 18420 14943 18472 14952
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 17592 14832 17644 14884
rect 2872 14764 2924 14816
rect 3884 14764 3936 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 14740 14764 14792 14816
rect 18052 14764 18104 14816
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 19892 15104 19944 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 24492 15104 24544 15156
rect 25044 15104 25096 15156
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 20904 15036 20956 15088
rect 22836 15011 22888 15020
rect 22836 14977 22845 15011
rect 22845 14977 22879 15011
rect 22879 14977 22888 15011
rect 24032 15036 24084 15088
rect 22836 14968 22888 14977
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 19248 14943 19300 14952
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 24492 14900 24544 14952
rect 25044 14900 25096 14952
rect 25872 14900 25924 14952
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 18880 14807 18932 14816
rect 18880 14773 18889 14807
rect 18889 14773 18923 14807
rect 18923 14773 18932 14807
rect 18880 14764 18932 14773
rect 19156 14764 19208 14816
rect 22468 14832 22520 14884
rect 23204 14832 23256 14884
rect 20720 14764 20772 14816
rect 22744 14807 22796 14816
rect 22744 14773 22753 14807
rect 22753 14773 22787 14807
rect 22787 14773 22796 14807
rect 22744 14764 22796 14773
rect 24124 14832 24176 14884
rect 24584 14832 24636 14884
rect 24216 14764 24268 14816
rect 4169 14662 4221 14714
rect 4233 14662 4285 14714
rect 4297 14662 4349 14714
rect 4361 14662 4413 14714
rect 4425 14662 4477 14714
rect 10608 14662 10660 14714
rect 10672 14662 10724 14714
rect 10736 14662 10788 14714
rect 10800 14662 10852 14714
rect 10864 14662 10916 14714
rect 17047 14662 17099 14714
rect 17111 14662 17163 14714
rect 17175 14662 17227 14714
rect 17239 14662 17291 14714
rect 17303 14662 17355 14714
rect 23486 14662 23538 14714
rect 23550 14662 23602 14714
rect 23614 14662 23666 14714
rect 23678 14662 23730 14714
rect 23742 14662 23794 14714
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 15108 14560 15160 14612
rect 15936 14560 15988 14612
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 17684 14603 17736 14612
rect 3332 14492 3384 14544
rect 3700 14492 3752 14544
rect 10232 14492 10284 14544
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 3424 14424 3476 14476
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5264 14288 5316 14340
rect 7196 14356 7248 14408
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 2780 14220 2832 14229
rect 3332 14220 3384 14272
rect 3976 14220 4028 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 6644 14220 6696 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 7656 14288 7708 14340
rect 7932 14356 7984 14408
rect 8484 14424 8536 14476
rect 8852 14356 8904 14408
rect 9404 14399 9456 14408
rect 9404 14365 9413 14399
rect 9413 14365 9447 14399
rect 9447 14365 9456 14399
rect 9404 14356 9456 14365
rect 14556 14424 14608 14476
rect 17684 14569 17693 14603
rect 17693 14569 17727 14603
rect 17727 14569 17736 14603
rect 17684 14560 17736 14569
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 13636 14356 13688 14408
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 14924 14356 14976 14408
rect 16580 14356 16632 14408
rect 16856 14356 16908 14408
rect 17408 14356 17460 14408
rect 18052 14424 18104 14476
rect 18420 14492 18472 14544
rect 18880 14560 18932 14612
rect 19524 14560 19576 14612
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 19064 14492 19116 14544
rect 19892 14492 19944 14544
rect 20628 14560 20680 14612
rect 24860 14560 24912 14612
rect 18972 14424 19024 14476
rect 19800 14424 19852 14476
rect 20720 14424 20772 14476
rect 23940 14424 23992 14476
rect 8760 14288 8812 14340
rect 12256 14288 12308 14340
rect 15660 14288 15712 14340
rect 18328 14377 18380 14386
rect 18328 14343 18337 14377
rect 18337 14343 18371 14377
rect 18371 14343 18380 14377
rect 18328 14334 18380 14343
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8668 14220 8720 14272
rect 9772 14220 9824 14272
rect 11704 14220 11756 14272
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 15568 14263 15620 14272
rect 15568 14229 15577 14263
rect 15577 14229 15611 14263
rect 15611 14229 15620 14263
rect 15568 14220 15620 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 16672 14220 16724 14272
rect 17500 14263 17552 14272
rect 17500 14229 17509 14263
rect 17509 14229 17543 14263
rect 17543 14229 17552 14263
rect 17500 14220 17552 14229
rect 19064 14399 19116 14408
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 19156 14356 19208 14408
rect 18696 14288 18748 14340
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 22560 14399 22612 14408
rect 22560 14365 22569 14399
rect 22569 14365 22603 14399
rect 22603 14365 22612 14399
rect 22560 14356 22612 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 22928 14356 22980 14408
rect 23204 14356 23256 14408
rect 24216 14399 24268 14408
rect 24216 14365 24225 14399
rect 24225 14365 24259 14399
rect 24259 14365 24268 14399
rect 24216 14356 24268 14365
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 24124 14288 24176 14340
rect 18788 14220 18840 14272
rect 19432 14220 19484 14272
rect 22192 14220 22244 14272
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 23848 14220 23900 14272
rect 25044 14288 25096 14340
rect 25964 14263 26016 14272
rect 25964 14229 25973 14263
rect 25973 14229 26007 14263
rect 26007 14229 26016 14263
rect 25964 14220 26016 14229
rect 4829 14118 4881 14170
rect 4893 14118 4945 14170
rect 4957 14118 5009 14170
rect 5021 14118 5073 14170
rect 5085 14118 5137 14170
rect 11268 14118 11320 14170
rect 11332 14118 11384 14170
rect 11396 14118 11448 14170
rect 11460 14118 11512 14170
rect 11524 14118 11576 14170
rect 17707 14118 17759 14170
rect 17771 14118 17823 14170
rect 17835 14118 17887 14170
rect 17899 14118 17951 14170
rect 17963 14118 18015 14170
rect 24146 14118 24198 14170
rect 24210 14118 24262 14170
rect 24274 14118 24326 14170
rect 24338 14118 24390 14170
rect 24402 14118 24454 14170
rect 3700 14016 3752 14068
rect 4252 14016 4304 14068
rect 3148 13948 3200 14000
rect 6552 14016 6604 14068
rect 6920 14016 6972 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 8484 14016 8536 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 13636 14059 13688 14068
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 14556 14059 14608 14068
rect 14556 14025 14565 14059
rect 14565 14025 14599 14059
rect 14599 14025 14608 14059
rect 14556 14016 14608 14025
rect 14924 14016 14976 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 4068 13880 4120 13932
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 5172 13880 5224 13932
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 7104 13991 7156 14000
rect 7104 13957 7113 13991
rect 7113 13957 7147 13991
rect 7147 13957 7156 13991
rect 7104 13948 7156 13957
rect 7932 13948 7984 14000
rect 8208 13948 8260 14000
rect 7472 13880 7524 13932
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 3976 13744 4028 13796
rect 5540 13812 5592 13864
rect 7104 13812 7156 13864
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 8576 13880 8628 13932
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 10048 13991 10100 14000
rect 10048 13957 10057 13991
rect 10057 13957 10091 13991
rect 10091 13957 10100 13991
rect 10048 13948 10100 13957
rect 11612 13880 11664 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12072 13948 12124 14000
rect 13544 13948 13596 14000
rect 15016 13948 15068 14000
rect 18144 14016 18196 14068
rect 18696 14016 18748 14068
rect 22560 14016 22612 14068
rect 22652 14016 22704 14068
rect 24860 14059 24912 14068
rect 24860 14025 24869 14059
rect 24869 14025 24903 14059
rect 24903 14025 24912 14059
rect 24860 14016 24912 14025
rect 25320 14016 25372 14068
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 14924 13880 14976 13932
rect 18328 13948 18380 14000
rect 18604 13923 18656 13932
rect 4528 13787 4580 13796
rect 4528 13753 4537 13787
rect 4537 13753 4571 13787
rect 4571 13753 4580 13787
rect 4528 13744 4580 13753
rect 7564 13744 7616 13796
rect 8852 13812 8904 13864
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 9128 13744 9180 13796
rect 13176 13744 13228 13796
rect 15016 13812 15068 13864
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 17500 13812 17552 13864
rect 18328 13812 18380 13864
rect 1676 13676 1728 13728
rect 2780 13676 2832 13728
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 4712 13676 4764 13728
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 6460 13719 6512 13728
rect 6460 13685 6469 13719
rect 6469 13685 6503 13719
rect 6503 13685 6512 13719
rect 6460 13676 6512 13685
rect 7840 13676 7892 13728
rect 8852 13676 8904 13728
rect 10048 13676 10100 13728
rect 11060 13676 11112 13728
rect 11152 13676 11204 13728
rect 14832 13676 14884 13728
rect 18052 13744 18104 13796
rect 19800 13812 19852 13864
rect 22100 13812 22152 13864
rect 22744 13880 22796 13932
rect 24492 13948 24544 14000
rect 23020 13880 23072 13932
rect 23296 13923 23348 13932
rect 23296 13889 23305 13923
rect 23305 13889 23339 13923
rect 23339 13889 23348 13923
rect 23296 13880 23348 13889
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 23756 13880 23808 13932
rect 25964 13880 26016 13932
rect 22928 13812 22980 13864
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 23020 13744 23072 13796
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 16948 13676 17000 13728
rect 18880 13676 18932 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 4169 13574 4221 13626
rect 4233 13574 4285 13626
rect 4297 13574 4349 13626
rect 4361 13574 4413 13626
rect 4425 13574 4477 13626
rect 10608 13574 10660 13626
rect 10672 13574 10724 13626
rect 10736 13574 10788 13626
rect 10800 13574 10852 13626
rect 10864 13574 10916 13626
rect 17047 13574 17099 13626
rect 17111 13574 17163 13626
rect 17175 13574 17227 13626
rect 17239 13574 17291 13626
rect 17303 13574 17355 13626
rect 23486 13574 23538 13626
rect 23550 13574 23602 13626
rect 23614 13574 23666 13626
rect 23678 13574 23730 13626
rect 23742 13574 23794 13626
rect 3240 13515 3292 13524
rect 3240 13481 3249 13515
rect 3249 13481 3283 13515
rect 3283 13481 3292 13515
rect 3240 13472 3292 13481
rect 3976 13515 4028 13524
rect 3976 13481 3985 13515
rect 3985 13481 4019 13515
rect 4019 13481 4028 13515
rect 3976 13472 4028 13481
rect 4160 13515 4212 13524
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 4988 13472 5040 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 7104 13472 7156 13524
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 4344 13404 4396 13456
rect 4160 13336 4212 13388
rect 1676 13268 1728 13320
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2688 13268 2740 13320
rect 3240 13268 3292 13320
rect 3884 13200 3936 13252
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 5632 13336 5684 13388
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6460 13268 6512 13320
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 8116 13336 8168 13388
rect 8576 13404 8628 13456
rect 8852 13404 8904 13456
rect 12808 13472 12860 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 15016 13472 15068 13524
rect 15384 13472 15436 13524
rect 18880 13472 18932 13524
rect 5448 13200 5500 13252
rect 7932 13268 7984 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 11612 13336 11664 13388
rect 12072 13336 12124 13388
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 17500 13404 17552 13456
rect 22100 13472 22152 13524
rect 22836 13472 22888 13524
rect 24124 13472 24176 13524
rect 8300 13200 8352 13252
rect 7380 13132 7432 13184
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 8852 13268 8904 13320
rect 10048 13311 10100 13320
rect 10048 13277 10066 13311
rect 10066 13277 10100 13311
rect 10048 13268 10100 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 12348 13268 12400 13320
rect 13268 13268 13320 13320
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 16120 13336 16172 13388
rect 18052 13336 18104 13388
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 19248 13336 19300 13388
rect 20628 13336 20680 13388
rect 23204 13404 23256 13456
rect 23848 13447 23900 13456
rect 23848 13413 23857 13447
rect 23857 13413 23891 13447
rect 23891 13413 23900 13447
rect 23848 13404 23900 13413
rect 23940 13404 23992 13456
rect 23020 13336 23072 13388
rect 23296 13336 23348 13388
rect 18144 13268 18196 13320
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 23388 13268 23440 13320
rect 24584 13336 24636 13388
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 11152 13200 11204 13252
rect 15752 13200 15804 13252
rect 16948 13200 17000 13252
rect 15016 13132 15068 13184
rect 15292 13132 15344 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 16120 13132 16172 13184
rect 18144 13132 18196 13184
rect 20076 13200 20128 13252
rect 24952 13243 25004 13252
rect 24952 13209 24986 13243
rect 24986 13209 25004 13243
rect 24952 13200 25004 13209
rect 26240 13132 26292 13184
rect 4829 13030 4881 13082
rect 4893 13030 4945 13082
rect 4957 13030 5009 13082
rect 5021 13030 5073 13082
rect 5085 13030 5137 13082
rect 11268 13030 11320 13082
rect 11332 13030 11384 13082
rect 11396 13030 11448 13082
rect 11460 13030 11512 13082
rect 11524 13030 11576 13082
rect 17707 13030 17759 13082
rect 17771 13030 17823 13082
rect 17835 13030 17887 13082
rect 17899 13030 17951 13082
rect 17963 13030 18015 13082
rect 24146 13030 24198 13082
rect 24210 13030 24262 13082
rect 24274 13030 24326 13082
rect 24338 13030 24390 13082
rect 24402 13030 24454 13082
rect 3424 12928 3476 12980
rect 3792 12928 3844 12980
rect 3884 12928 3936 12980
rect 3976 12903 4028 12912
rect 3976 12869 3985 12903
rect 3985 12869 4019 12903
rect 4019 12869 4028 12903
rect 3976 12860 4028 12869
rect 4344 12860 4396 12912
rect 5264 12903 5316 12912
rect 5264 12869 5273 12903
rect 5273 12869 5307 12903
rect 5307 12869 5316 12903
rect 5264 12860 5316 12869
rect 7564 12928 7616 12980
rect 7932 12928 7984 12980
rect 8576 12928 8628 12980
rect 9404 12860 9456 12912
rect 11428 12928 11480 12980
rect 11704 12928 11756 12980
rect 12164 12928 12216 12980
rect 13268 12928 13320 12980
rect 15568 12928 15620 12980
rect 15752 12928 15804 12980
rect 17500 12928 17552 12980
rect 20076 12928 20128 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 23940 12928 23992 12980
rect 24676 12928 24728 12980
rect 24952 12928 25004 12980
rect 11060 12903 11112 12912
rect 11060 12869 11069 12903
rect 11069 12869 11103 12903
rect 11103 12869 11112 12903
rect 11060 12860 11112 12869
rect 12072 12860 12124 12912
rect 13452 12860 13504 12912
rect 15476 12860 15528 12912
rect 15936 12860 15988 12912
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 3332 12792 3384 12844
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 4528 12792 4580 12844
rect 4620 12792 4672 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 5448 12792 5500 12844
rect 7104 12792 7156 12844
rect 7840 12792 7892 12844
rect 8024 12792 8076 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 11612 12792 11664 12844
rect 12256 12792 12308 12844
rect 13176 12792 13228 12844
rect 15292 12792 15344 12844
rect 5632 12724 5684 12776
rect 8116 12724 8168 12776
rect 8760 12724 8812 12776
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 4620 12699 4672 12708
rect 4620 12665 4629 12699
rect 4629 12665 4663 12699
rect 4663 12665 4672 12699
rect 4620 12656 4672 12665
rect 5172 12656 5224 12708
rect 9036 12699 9088 12708
rect 9036 12665 9045 12699
rect 9045 12665 9079 12699
rect 9079 12665 9088 12699
rect 9036 12656 9088 12665
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 13268 12656 13320 12708
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 18696 12860 18748 12912
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 19064 12792 19116 12844
rect 3976 12588 4028 12640
rect 4436 12588 4488 12640
rect 9128 12588 9180 12640
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 15384 12588 15436 12640
rect 15752 12656 15804 12708
rect 18144 12724 18196 12776
rect 20812 12792 20864 12844
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 19984 12724 20036 12776
rect 20628 12767 20680 12776
rect 20628 12733 20637 12767
rect 20637 12733 20671 12767
rect 20671 12733 20680 12767
rect 20628 12724 20680 12733
rect 24860 12792 24912 12844
rect 25044 12835 25096 12844
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 25320 12835 25372 12844
rect 25320 12801 25329 12835
rect 25329 12801 25363 12835
rect 25363 12801 25372 12835
rect 25320 12792 25372 12801
rect 26240 12724 26292 12776
rect 20812 12656 20864 12708
rect 20996 12656 21048 12708
rect 16212 12588 16264 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 4169 12486 4221 12538
rect 4233 12486 4285 12538
rect 4297 12486 4349 12538
rect 4361 12486 4413 12538
rect 4425 12486 4477 12538
rect 10608 12486 10660 12538
rect 10672 12486 10724 12538
rect 10736 12486 10788 12538
rect 10800 12486 10852 12538
rect 10864 12486 10916 12538
rect 17047 12486 17099 12538
rect 17111 12486 17163 12538
rect 17175 12486 17227 12538
rect 17239 12486 17291 12538
rect 17303 12486 17355 12538
rect 23486 12486 23538 12538
rect 23550 12486 23602 12538
rect 23614 12486 23666 12538
rect 23678 12486 23730 12538
rect 23742 12486 23794 12538
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 4528 12384 4580 12436
rect 4620 12384 4672 12436
rect 8484 12384 8536 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12808 12384 12860 12436
rect 16948 12384 17000 12436
rect 20904 12384 20956 12436
rect 21640 12384 21692 12436
rect 2688 12316 2740 12368
rect 5172 12316 5224 12368
rect 5816 12316 5868 12368
rect 8392 12316 8444 12368
rect 21364 12316 21416 12368
rect 22008 12384 22060 12436
rect 22836 12427 22888 12436
rect 22836 12393 22845 12427
rect 22845 12393 22879 12427
rect 22879 12393 22888 12427
rect 22836 12384 22888 12393
rect 23388 12316 23440 12368
rect 3424 12248 3476 12300
rect 4160 12248 4212 12300
rect 7380 12248 7432 12300
rect 15384 12248 15436 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 17592 12248 17644 12300
rect 19064 12248 19116 12300
rect 2044 12180 2096 12232
rect 2320 12180 2372 12232
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 7656 12180 7708 12232
rect 8300 12180 8352 12232
rect 11796 12180 11848 12232
rect 12348 12180 12400 12232
rect 14648 12180 14700 12232
rect 18052 12180 18104 12232
rect 18788 12180 18840 12232
rect 9588 12112 9640 12164
rect 16764 12112 16816 12164
rect 19064 12112 19116 12164
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 20812 12248 20864 12300
rect 23020 12248 23072 12300
rect 21824 12180 21876 12232
rect 23112 12223 23164 12232
rect 23112 12189 23121 12223
rect 23121 12189 23155 12223
rect 23155 12189 23164 12223
rect 23112 12180 23164 12189
rect 19432 12112 19484 12164
rect 19524 12155 19576 12164
rect 19524 12121 19533 12155
rect 19533 12121 19567 12155
rect 19567 12121 19576 12155
rect 19524 12112 19576 12121
rect 20076 12112 20128 12164
rect 21456 12155 21508 12164
rect 21456 12121 21465 12155
rect 21465 12121 21499 12155
rect 21499 12121 21508 12155
rect 21456 12112 21508 12121
rect 17316 12044 17368 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 18236 12044 18288 12096
rect 18880 12044 18932 12096
rect 22652 12087 22704 12096
rect 22652 12053 22661 12087
rect 22661 12053 22695 12087
rect 22695 12053 22704 12087
rect 22652 12044 22704 12053
rect 4829 11942 4881 11994
rect 4893 11942 4945 11994
rect 4957 11942 5009 11994
rect 5021 11942 5073 11994
rect 5085 11942 5137 11994
rect 11268 11942 11320 11994
rect 11332 11942 11384 11994
rect 11396 11942 11448 11994
rect 11460 11942 11512 11994
rect 11524 11942 11576 11994
rect 17707 11942 17759 11994
rect 17771 11942 17823 11994
rect 17835 11942 17887 11994
rect 17899 11942 17951 11994
rect 17963 11942 18015 11994
rect 24146 11942 24198 11994
rect 24210 11942 24262 11994
rect 24274 11942 24326 11994
rect 24338 11942 24390 11994
rect 24402 11942 24454 11994
rect 14464 11840 14516 11892
rect 15292 11840 15344 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 15936 11772 15988 11824
rect 16120 11772 16172 11824
rect 18052 11840 18104 11892
rect 18880 11772 18932 11824
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 20904 11840 20956 11892
rect 21640 11772 21692 11824
rect 21732 11772 21784 11824
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 19432 11704 19484 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 22008 11704 22060 11756
rect 22376 11772 22428 11824
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22468 11704 22520 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 13728 11636 13780 11688
rect 12348 11500 12400 11552
rect 14556 11636 14608 11688
rect 16488 11679 16540 11688
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 22928 11679 22980 11688
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 25780 11704 25832 11756
rect 26516 11747 26568 11756
rect 26516 11713 26525 11747
rect 26525 11713 26559 11747
rect 26559 11713 26568 11747
rect 26516 11704 26568 11713
rect 16672 11500 16724 11552
rect 21456 11568 21508 11620
rect 21824 11568 21876 11620
rect 21732 11500 21784 11552
rect 23940 11500 23992 11552
rect 26332 11543 26384 11552
rect 26332 11509 26341 11543
rect 26341 11509 26375 11543
rect 26375 11509 26384 11543
rect 26332 11500 26384 11509
rect 4169 11398 4221 11450
rect 4233 11398 4285 11450
rect 4297 11398 4349 11450
rect 4361 11398 4413 11450
rect 4425 11398 4477 11450
rect 10608 11398 10660 11450
rect 10672 11398 10724 11450
rect 10736 11398 10788 11450
rect 10800 11398 10852 11450
rect 10864 11398 10916 11450
rect 17047 11398 17099 11450
rect 17111 11398 17163 11450
rect 17175 11398 17227 11450
rect 17239 11398 17291 11450
rect 17303 11398 17355 11450
rect 23486 11398 23538 11450
rect 23550 11398 23602 11450
rect 23614 11398 23666 11450
rect 23678 11398 23730 11450
rect 23742 11398 23794 11450
rect 9220 11296 9272 11348
rect 3516 11228 3568 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4068 11160 4120 11212
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 5448 11160 5500 11212
rect 8576 11160 8628 11212
rect 2964 11067 3016 11076
rect 2964 11033 2973 11067
rect 2973 11033 3007 11067
rect 3007 11033 3016 11067
rect 11152 11092 11204 11144
rect 15936 11296 15988 11348
rect 19524 11296 19576 11348
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22192 11296 22244 11348
rect 22744 11296 22796 11348
rect 22928 11339 22980 11348
rect 22928 11305 22937 11339
rect 22937 11305 22971 11339
rect 22971 11305 22980 11339
rect 22928 11296 22980 11305
rect 23204 11296 23256 11348
rect 16028 11228 16080 11280
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 15568 11160 15620 11212
rect 16488 11160 16540 11212
rect 19248 11203 19300 11212
rect 19248 11169 19257 11203
rect 19257 11169 19291 11203
rect 19291 11169 19300 11203
rect 19248 11160 19300 11169
rect 22192 11160 22244 11212
rect 23388 11228 23440 11280
rect 23940 11296 23992 11348
rect 2964 11024 3016 11033
rect 3884 11024 3936 11076
rect 5356 11024 5408 11076
rect 6460 11024 6512 11076
rect 11060 11024 11112 11076
rect 14556 11092 14608 11144
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 18420 11092 18472 11144
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 22468 11092 22520 11144
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 24584 11092 24636 11144
rect 25780 11092 25832 11144
rect 13084 11024 13136 11076
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 19616 11024 19668 11076
rect 23020 11024 23072 11076
rect 23204 11067 23256 11076
rect 23204 11033 23213 11067
rect 23213 11033 23247 11067
rect 23247 11033 23256 11067
rect 23204 11024 23256 11033
rect 3424 10999 3476 11008
rect 3424 10965 3433 10999
rect 3433 10965 3467 10999
rect 3467 10965 3476 10999
rect 3424 10956 3476 10965
rect 6368 10956 6420 11008
rect 6736 10956 6788 11008
rect 8760 10956 8812 11008
rect 9956 10956 10008 11008
rect 13636 10956 13688 11008
rect 14188 10999 14240 11008
rect 14188 10965 14197 10999
rect 14197 10965 14231 10999
rect 14231 10965 14240 10999
rect 14188 10956 14240 10965
rect 24860 10999 24912 11008
rect 24860 10965 24869 10999
rect 24869 10965 24903 10999
rect 24903 10965 24912 10999
rect 24860 10956 24912 10965
rect 4829 10854 4881 10906
rect 4893 10854 4945 10906
rect 4957 10854 5009 10906
rect 5021 10854 5073 10906
rect 5085 10854 5137 10906
rect 11268 10854 11320 10906
rect 11332 10854 11384 10906
rect 11396 10854 11448 10906
rect 11460 10854 11512 10906
rect 11524 10854 11576 10906
rect 17707 10854 17759 10906
rect 17771 10854 17823 10906
rect 17835 10854 17887 10906
rect 17899 10854 17951 10906
rect 17963 10854 18015 10906
rect 24146 10854 24198 10906
rect 24210 10854 24262 10906
rect 24274 10854 24326 10906
rect 24338 10854 24390 10906
rect 24402 10854 24454 10906
rect 4252 10752 4304 10804
rect 5264 10752 5316 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 1860 10684 1912 10736
rect 3424 10684 3476 10736
rect 5540 10727 5592 10736
rect 5540 10693 5549 10727
rect 5549 10693 5583 10727
rect 5583 10693 5592 10727
rect 5540 10684 5592 10693
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 3976 10616 4028 10668
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 4896 10616 4948 10668
rect 4620 10548 4672 10600
rect 5264 10616 5316 10668
rect 5908 10616 5960 10668
rect 6368 10616 6420 10668
rect 8024 10752 8076 10804
rect 8116 10752 8168 10804
rect 8668 10752 8720 10804
rect 8760 10752 8812 10804
rect 6828 10684 6880 10736
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 7472 10616 7524 10668
rect 9404 10684 9456 10736
rect 11152 10752 11204 10804
rect 13084 10752 13136 10804
rect 15660 10752 15712 10804
rect 19616 10795 19668 10804
rect 19616 10761 19625 10795
rect 19625 10761 19659 10795
rect 19659 10761 19668 10795
rect 19616 10752 19668 10761
rect 22560 10752 22612 10804
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8576 10616 8628 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 10416 10616 10468 10668
rect 11152 10616 11204 10668
rect 11796 10616 11848 10668
rect 14464 10684 14516 10736
rect 21824 10727 21876 10736
rect 21824 10693 21833 10727
rect 21833 10693 21867 10727
rect 21867 10693 21876 10727
rect 21824 10684 21876 10693
rect 6920 10548 6972 10600
rect 8944 10548 8996 10600
rect 9036 10591 9088 10600
rect 9036 10557 9045 10591
rect 9045 10557 9079 10591
rect 9079 10557 9088 10591
rect 9036 10548 9088 10557
rect 4068 10480 4120 10532
rect 4712 10480 4764 10532
rect 5080 10480 5132 10532
rect 3700 10412 3752 10464
rect 4620 10455 4672 10464
rect 4620 10421 4629 10455
rect 4629 10421 4663 10455
rect 4663 10421 4672 10455
rect 4620 10412 4672 10421
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 5632 10480 5684 10532
rect 8208 10480 8260 10532
rect 7840 10412 7892 10464
rect 8576 10480 8628 10532
rect 8760 10480 8812 10532
rect 9404 10548 9456 10600
rect 11704 10548 11756 10600
rect 12072 10591 12124 10600
rect 12072 10557 12081 10591
rect 12081 10557 12115 10591
rect 12115 10557 12124 10591
rect 12072 10548 12124 10557
rect 15292 10616 15344 10668
rect 19432 10616 19484 10668
rect 22100 10616 22152 10668
rect 22928 10659 22980 10668
rect 14464 10548 14516 10600
rect 14740 10591 14792 10600
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 8668 10412 8720 10464
rect 9496 10412 9548 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 22192 10455 22244 10464
rect 22192 10421 22201 10455
rect 22201 10421 22235 10455
rect 22235 10421 22244 10455
rect 22192 10412 22244 10421
rect 22284 10455 22336 10464
rect 22284 10421 22293 10455
rect 22293 10421 22327 10455
rect 22327 10421 22336 10455
rect 22284 10412 22336 10421
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 24860 10752 24912 10804
rect 25780 10795 25832 10804
rect 25780 10761 25789 10795
rect 25789 10761 25823 10795
rect 25823 10761 25832 10795
rect 25780 10752 25832 10761
rect 22744 10412 22796 10464
rect 24032 10412 24084 10464
rect 24492 10616 24544 10668
rect 25044 10412 25096 10464
rect 4169 10310 4221 10362
rect 4233 10310 4285 10362
rect 4297 10310 4349 10362
rect 4361 10310 4413 10362
rect 4425 10310 4477 10362
rect 10608 10310 10660 10362
rect 10672 10310 10724 10362
rect 10736 10310 10788 10362
rect 10800 10310 10852 10362
rect 10864 10310 10916 10362
rect 17047 10310 17099 10362
rect 17111 10310 17163 10362
rect 17175 10310 17227 10362
rect 17239 10310 17291 10362
rect 17303 10310 17355 10362
rect 23486 10310 23538 10362
rect 23550 10310 23602 10362
rect 23614 10310 23666 10362
rect 23678 10310 23730 10362
rect 23742 10310 23794 10362
rect 4068 10208 4120 10260
rect 5080 10208 5132 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 4620 10140 4672 10192
rect 1860 10072 1912 10124
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5264 10072 5316 10124
rect 7748 10208 7800 10260
rect 8760 10208 8812 10260
rect 9496 10208 9548 10260
rect 12072 10208 12124 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 21824 10208 21876 10260
rect 5816 10140 5868 10192
rect 6828 10140 6880 10192
rect 8484 10140 8536 10192
rect 8576 10140 8628 10192
rect 13728 10183 13780 10192
rect 13728 10149 13737 10183
rect 13737 10149 13771 10183
rect 13771 10149 13780 10183
rect 13728 10140 13780 10149
rect 14464 10140 14516 10192
rect 22192 10208 22244 10260
rect 22376 10208 22428 10260
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 4804 10004 4856 10056
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 2872 9936 2924 9988
rect 4252 9979 4304 9988
rect 4252 9945 4261 9979
rect 4261 9945 4295 9979
rect 4295 9945 4304 9979
rect 4252 9936 4304 9945
rect 4344 9979 4396 9988
rect 4344 9945 4353 9979
rect 4353 9945 4387 9979
rect 4387 9945 4396 9979
rect 4344 9936 4396 9945
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6368 9936 6420 9988
rect 6460 9979 6512 9988
rect 6460 9945 6469 9979
rect 6469 9945 6503 9979
rect 6503 9945 6512 9979
rect 6460 9936 6512 9945
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7472 10004 7524 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 7840 10004 7892 10056
rect 9036 10072 9088 10124
rect 10324 10072 10376 10124
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 8208 10004 8260 10056
rect 7564 9936 7616 9988
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9312 10004 9364 10056
rect 9496 10004 9548 10056
rect 13636 10004 13688 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15200 10004 15252 10056
rect 19432 10004 19484 10056
rect 24492 10072 24544 10124
rect 4988 9868 5040 9920
rect 6000 9868 6052 9920
rect 7840 9868 7892 9920
rect 7932 9868 7984 9920
rect 9956 9979 10008 9988
rect 9956 9945 9965 9979
rect 9965 9945 9999 9979
rect 9999 9945 10008 9979
rect 9956 9936 10008 9945
rect 11244 9936 11296 9988
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8944 9868 8996 9920
rect 11888 9979 11940 9988
rect 11888 9945 11897 9979
rect 11897 9945 11931 9979
rect 11931 9945 11940 9979
rect 11888 9936 11940 9945
rect 12440 9936 12492 9988
rect 21272 9936 21324 9988
rect 21364 9936 21416 9988
rect 21916 9936 21968 9988
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 25320 10004 25372 10056
rect 24768 9936 24820 9988
rect 12900 9868 12952 9920
rect 22100 9911 22152 9920
rect 22100 9877 22109 9911
rect 22109 9877 22143 9911
rect 22143 9877 22152 9911
rect 22100 9868 22152 9877
rect 23020 9868 23072 9920
rect 25136 9868 25188 9920
rect 26056 9911 26108 9920
rect 26056 9877 26065 9911
rect 26065 9877 26099 9911
rect 26099 9877 26108 9911
rect 26056 9868 26108 9877
rect 4829 9766 4881 9818
rect 4893 9766 4945 9818
rect 4957 9766 5009 9818
rect 5021 9766 5073 9818
rect 5085 9766 5137 9818
rect 11268 9766 11320 9818
rect 11332 9766 11384 9818
rect 11396 9766 11448 9818
rect 11460 9766 11512 9818
rect 11524 9766 11576 9818
rect 17707 9766 17759 9818
rect 17771 9766 17823 9818
rect 17835 9766 17887 9818
rect 17899 9766 17951 9818
rect 17963 9766 18015 9818
rect 24146 9766 24198 9818
rect 24210 9766 24262 9818
rect 24274 9766 24326 9818
rect 24338 9766 24390 9818
rect 24402 9766 24454 9818
rect 4252 9664 4304 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 6368 9664 6420 9716
rect 8024 9664 8076 9716
rect 3700 9596 3752 9648
rect 1860 9528 1912 9580
rect 4528 9596 4580 9648
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5172 9528 5224 9580
rect 5816 9528 5868 9580
rect 6184 9639 6236 9648
rect 6184 9605 6193 9639
rect 6193 9605 6227 9639
rect 6227 9605 6236 9639
rect 6184 9596 6236 9605
rect 4344 9460 4396 9512
rect 6000 9460 6052 9512
rect 6460 9528 6512 9580
rect 6920 9596 6972 9648
rect 7840 9639 7892 9648
rect 7840 9605 7849 9639
rect 7849 9605 7883 9639
rect 7883 9605 7892 9639
rect 7840 9596 7892 9605
rect 7932 9639 7984 9648
rect 7932 9605 7941 9639
rect 7941 9605 7975 9639
rect 7975 9605 7984 9639
rect 7932 9596 7984 9605
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 7472 9528 7524 9580
rect 7748 9528 7800 9580
rect 8392 9528 8444 9580
rect 9312 9596 9364 9648
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 8576 9528 8628 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 8944 9528 8996 9580
rect 21272 9707 21324 9716
rect 21272 9673 21281 9707
rect 21281 9673 21315 9707
rect 21315 9673 21324 9707
rect 21272 9664 21324 9673
rect 21916 9707 21968 9716
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 22100 9664 22152 9716
rect 24032 9707 24084 9716
rect 24032 9673 24041 9707
rect 24041 9673 24075 9707
rect 24075 9673 24084 9707
rect 24032 9664 24084 9673
rect 25320 9707 25372 9716
rect 25320 9673 25329 9707
rect 25329 9673 25363 9707
rect 25363 9673 25372 9707
rect 25320 9664 25372 9673
rect 10416 9596 10468 9648
rect 12440 9596 12492 9648
rect 15568 9596 15620 9648
rect 16672 9596 16724 9648
rect 11152 9528 11204 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 7564 9460 7616 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 19432 9528 19484 9580
rect 22928 9596 22980 9648
rect 21732 9528 21784 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 22744 9503 22796 9512
rect 22744 9469 22753 9503
rect 22753 9469 22787 9503
rect 22787 9469 22796 9503
rect 22744 9460 22796 9469
rect 23204 9596 23256 9648
rect 25044 9596 25096 9648
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 24768 9528 24820 9580
rect 23388 9460 23440 9512
rect 24584 9460 24636 9512
rect 26056 9528 26108 9580
rect 3976 9324 4028 9376
rect 5172 9324 5224 9376
rect 5264 9324 5316 9376
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 5908 9324 5960 9376
rect 6092 9324 6144 9376
rect 7012 9324 7064 9376
rect 11888 9324 11940 9376
rect 12808 9324 12860 9376
rect 13820 9324 13872 9376
rect 15752 9324 15804 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 22192 9367 22244 9376
rect 22192 9333 22201 9367
rect 22201 9333 22235 9367
rect 22235 9333 22244 9367
rect 22192 9324 22244 9333
rect 23204 9367 23256 9376
rect 23204 9333 23213 9367
rect 23213 9333 23247 9367
rect 23247 9333 23256 9367
rect 23204 9324 23256 9333
rect 23940 9392 23992 9444
rect 24584 9324 24636 9376
rect 25136 9367 25188 9376
rect 25136 9333 25145 9367
rect 25145 9333 25179 9367
rect 25179 9333 25188 9367
rect 25136 9324 25188 9333
rect 4169 9222 4221 9274
rect 4233 9222 4285 9274
rect 4297 9222 4349 9274
rect 4361 9222 4413 9274
rect 4425 9222 4477 9274
rect 10608 9222 10660 9274
rect 10672 9222 10724 9274
rect 10736 9222 10788 9274
rect 10800 9222 10852 9274
rect 10864 9222 10916 9274
rect 17047 9222 17099 9274
rect 17111 9222 17163 9274
rect 17175 9222 17227 9274
rect 17239 9222 17291 9274
rect 17303 9222 17355 9274
rect 23486 9222 23538 9274
rect 23550 9222 23602 9274
rect 23614 9222 23666 9274
rect 23678 9222 23730 9274
rect 23742 9222 23794 9274
rect 2872 9120 2924 9172
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 7104 9120 7156 9172
rect 11060 9120 11112 9172
rect 4620 9052 4672 9104
rect 5448 9052 5500 9104
rect 6184 9052 6236 9104
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 5908 8984 5960 9036
rect 8668 8984 8720 9036
rect 12808 9052 12860 9104
rect 13084 9120 13136 9172
rect 13728 9120 13780 9172
rect 14096 9120 14148 9172
rect 15568 9120 15620 9172
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 18144 9120 18196 9172
rect 18420 9120 18472 9172
rect 22192 9120 22244 9172
rect 23204 9120 23256 9172
rect 13636 9052 13688 9104
rect 940 8916 992 8968
rect 2964 8916 3016 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 10140 8848 10192 8900
rect 10784 8891 10836 8900
rect 10784 8857 10793 8891
rect 10793 8857 10827 8891
rect 10827 8857 10836 8891
rect 10784 8848 10836 8857
rect 11704 8848 11756 8900
rect 12900 8848 12952 8900
rect 13176 8891 13228 8900
rect 13176 8857 13185 8891
rect 13185 8857 13219 8891
rect 13219 8857 13228 8891
rect 13176 8848 13228 8857
rect 13268 8891 13320 8900
rect 13268 8857 13277 8891
rect 13277 8857 13311 8891
rect 13311 8857 13320 8891
rect 13268 8848 13320 8857
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 16028 8916 16080 8968
rect 15384 8848 15436 8900
rect 16764 8916 16816 8968
rect 17224 8916 17276 8968
rect 18052 8984 18104 9036
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 19248 9052 19300 9104
rect 19432 9052 19484 9104
rect 21824 8984 21876 9036
rect 23296 9052 23348 9104
rect 24032 9095 24084 9104
rect 24032 9061 24041 9095
rect 24041 9061 24075 9095
rect 24075 9061 24084 9095
rect 24032 9052 24084 9061
rect 2136 8780 2188 8832
rect 8576 8780 8628 8832
rect 12072 8780 12124 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 15108 8780 15160 8832
rect 18144 8780 18196 8832
rect 18420 8891 18472 8900
rect 18420 8857 18429 8891
rect 18429 8857 18463 8891
rect 18463 8857 18472 8891
rect 18420 8848 18472 8857
rect 18328 8780 18380 8832
rect 18512 8780 18564 8832
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 20352 8848 20404 8900
rect 24492 8984 24544 9036
rect 21272 8848 21324 8900
rect 26332 8916 26384 8968
rect 22100 8848 22152 8900
rect 22468 8848 22520 8900
rect 19340 8823 19392 8832
rect 19340 8789 19349 8823
rect 19349 8789 19383 8823
rect 19383 8789 19392 8823
rect 19340 8780 19392 8789
rect 20536 8823 20588 8832
rect 20536 8789 20545 8823
rect 20545 8789 20579 8823
rect 20579 8789 20588 8823
rect 20536 8780 20588 8789
rect 21732 8823 21784 8832
rect 21732 8789 21741 8823
rect 21741 8789 21775 8823
rect 21775 8789 21784 8823
rect 21732 8780 21784 8789
rect 22652 8780 22704 8832
rect 23388 8823 23440 8832
rect 23388 8789 23397 8823
rect 23397 8789 23431 8823
rect 23431 8789 23440 8823
rect 23388 8780 23440 8789
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 4829 8678 4881 8730
rect 4893 8678 4945 8730
rect 4957 8678 5009 8730
rect 5021 8678 5073 8730
rect 5085 8678 5137 8730
rect 11268 8678 11320 8730
rect 11332 8678 11384 8730
rect 11396 8678 11448 8730
rect 11460 8678 11512 8730
rect 11524 8678 11576 8730
rect 17707 8678 17759 8730
rect 17771 8678 17823 8730
rect 17835 8678 17887 8730
rect 17899 8678 17951 8730
rect 17963 8678 18015 8730
rect 24146 8678 24198 8730
rect 24210 8678 24262 8730
rect 24274 8678 24326 8730
rect 24338 8678 24390 8730
rect 24402 8678 24454 8730
rect 6184 8576 6236 8628
rect 13176 8576 13228 8628
rect 13728 8576 13780 8628
rect 14188 8576 14240 8628
rect 15016 8576 15068 8628
rect 17316 8576 17368 8628
rect 9128 8508 9180 8560
rect 12808 8508 12860 8560
rect 13452 8508 13504 8560
rect 14464 8508 14516 8560
rect 15752 8508 15804 8560
rect 18328 8576 18380 8628
rect 19524 8576 19576 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 5540 8440 5592 8492
rect 9036 8440 9088 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 8392 8304 8444 8356
rect 12900 8347 12952 8356
rect 12900 8313 12909 8347
rect 12909 8313 12943 8347
rect 12943 8313 12952 8347
rect 12900 8304 12952 8313
rect 13636 8440 13688 8492
rect 15292 8440 15344 8492
rect 17132 8440 17184 8492
rect 14096 8372 14148 8424
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18512 8508 18564 8560
rect 20536 8508 20588 8560
rect 18328 8440 18380 8492
rect 18696 8440 18748 8492
rect 9772 8236 9824 8288
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 13912 8236 13964 8288
rect 15016 8304 15068 8356
rect 17224 8304 17276 8356
rect 18972 8372 19024 8424
rect 19064 8372 19116 8424
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 20720 8440 20772 8492
rect 21732 8440 21784 8492
rect 23664 8508 23716 8560
rect 23940 8576 23992 8628
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 24492 8440 24544 8492
rect 19800 8415 19852 8424
rect 19800 8381 19809 8415
rect 19809 8381 19843 8415
rect 19843 8381 19852 8415
rect 19800 8372 19852 8381
rect 17960 8304 18012 8356
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18696 8347 18748 8356
rect 14096 8236 14148 8288
rect 14832 8236 14884 8288
rect 18696 8313 18705 8347
rect 18705 8313 18739 8347
rect 18739 8313 18748 8347
rect 18696 8304 18748 8313
rect 18420 8236 18472 8288
rect 19984 8236 20036 8288
rect 21640 8236 21692 8288
rect 4169 8134 4221 8186
rect 4233 8134 4285 8186
rect 4297 8134 4349 8186
rect 4361 8134 4413 8186
rect 4425 8134 4477 8186
rect 10608 8134 10660 8186
rect 10672 8134 10724 8186
rect 10736 8134 10788 8186
rect 10800 8134 10852 8186
rect 10864 8134 10916 8186
rect 17047 8134 17099 8186
rect 17111 8134 17163 8186
rect 17175 8134 17227 8186
rect 17239 8134 17291 8186
rect 17303 8134 17355 8186
rect 23486 8134 23538 8186
rect 23550 8134 23602 8186
rect 23614 8134 23666 8186
rect 23678 8134 23730 8186
rect 23742 8134 23794 8186
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 11980 8032 12032 8084
rect 12992 8032 13044 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 13636 8032 13688 8084
rect 14096 8075 14148 8084
rect 14096 8041 14105 8075
rect 14105 8041 14139 8075
rect 14139 8041 14148 8075
rect 14096 8032 14148 8041
rect 10968 7964 11020 8016
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 5632 7896 5684 7948
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 4528 7828 4580 7880
rect 9588 7896 9640 7948
rect 12716 7964 12768 8016
rect 7196 7828 7248 7880
rect 8300 7828 8352 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 10140 7828 10192 7880
rect 13452 7896 13504 7948
rect 13728 7896 13780 7948
rect 3792 7692 3844 7744
rect 7472 7760 7524 7812
rect 8208 7760 8260 7812
rect 9772 7760 9824 7812
rect 10692 7760 10744 7812
rect 11060 7803 11112 7812
rect 11060 7769 11069 7803
rect 11069 7769 11103 7803
rect 11103 7769 11112 7803
rect 11060 7760 11112 7769
rect 11888 7828 11940 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 13084 7828 13136 7880
rect 13636 7828 13688 7880
rect 14648 7871 14700 7880
rect 14648 7837 14652 7871
rect 14652 7837 14686 7871
rect 14686 7837 14700 7871
rect 14648 7828 14700 7837
rect 15016 7871 15068 7880
rect 15016 7837 15024 7871
rect 15024 7837 15058 7871
rect 15058 7837 15068 7871
rect 15016 7828 15068 7837
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 15752 7871 15804 7880
rect 15752 7837 15760 7871
rect 15760 7837 15794 7871
rect 15794 7837 15804 7871
rect 15752 7828 15804 7837
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 19800 8075 19852 8084
rect 19800 8041 19809 8075
rect 19809 8041 19843 8075
rect 19843 8041 19852 8075
rect 19800 8032 19852 8041
rect 20352 8032 20404 8084
rect 19340 7964 19392 8016
rect 20812 7964 20864 8016
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 19892 7896 19944 7948
rect 20076 7939 20128 7948
rect 20076 7905 20085 7939
rect 20085 7905 20119 7939
rect 20119 7905 20128 7939
rect 20076 7896 20128 7905
rect 20444 7896 20496 7948
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 20628 7896 20680 7948
rect 20996 7828 21048 7880
rect 11704 7760 11756 7812
rect 14464 7760 14516 7812
rect 14740 7803 14792 7812
rect 14740 7769 14749 7803
rect 14749 7769 14783 7803
rect 14783 7769 14792 7803
rect 14740 7760 14792 7769
rect 14832 7803 14884 7812
rect 14832 7769 14841 7803
rect 14841 7769 14875 7803
rect 14875 7769 14884 7803
rect 14832 7760 14884 7769
rect 8024 7692 8076 7744
rect 8760 7692 8812 7744
rect 11612 7692 11664 7744
rect 12440 7692 12492 7744
rect 15108 7692 15160 7744
rect 15200 7735 15252 7744
rect 15200 7701 15209 7735
rect 15209 7701 15243 7735
rect 15243 7701 15252 7735
rect 15200 7692 15252 7701
rect 15476 7803 15528 7812
rect 15476 7769 15485 7803
rect 15485 7769 15519 7803
rect 15519 7769 15528 7803
rect 15476 7760 15528 7769
rect 19800 7760 19852 7812
rect 18144 7692 18196 7744
rect 19892 7692 19944 7744
rect 20628 7692 20680 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 4829 7590 4881 7642
rect 4893 7590 4945 7642
rect 4957 7590 5009 7642
rect 5021 7590 5073 7642
rect 5085 7590 5137 7642
rect 11268 7590 11320 7642
rect 11332 7590 11384 7642
rect 11396 7590 11448 7642
rect 11460 7590 11512 7642
rect 11524 7590 11576 7642
rect 17707 7590 17759 7642
rect 17771 7590 17823 7642
rect 17835 7590 17887 7642
rect 17899 7590 17951 7642
rect 17963 7590 18015 7642
rect 24146 7590 24198 7642
rect 24210 7590 24262 7642
rect 24274 7590 24326 7642
rect 24338 7590 24390 7642
rect 24402 7590 24454 7642
rect 4252 7488 4304 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 3516 7420 3568 7472
rect 5632 7463 5684 7472
rect 5632 7429 5641 7463
rect 5641 7429 5675 7463
rect 5675 7429 5684 7463
rect 5632 7420 5684 7429
rect 3884 7284 3936 7336
rect 3240 7216 3292 7268
rect 4620 7352 4672 7404
rect 5356 7352 5408 7404
rect 5172 7284 5224 7336
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 8024 7420 8076 7472
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 12716 7488 12768 7540
rect 13728 7488 13780 7540
rect 14188 7488 14240 7540
rect 14648 7488 14700 7540
rect 16948 7488 17000 7540
rect 18788 7488 18840 7540
rect 19432 7488 19484 7540
rect 19800 7488 19852 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8944 7352 8996 7404
rect 8208 7284 8260 7336
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 7288 7216 7340 7268
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 10048 7284 10100 7336
rect 10140 7327 10192 7336
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 8668 7216 8720 7268
rect 10600 7284 10652 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 4804 7148 4856 7200
rect 5908 7148 5960 7200
rect 9128 7148 9180 7200
rect 9772 7148 9824 7200
rect 11152 7148 11204 7200
rect 13452 7420 13504 7472
rect 11796 7352 11848 7404
rect 13636 7352 13688 7404
rect 14004 7420 14056 7472
rect 19984 7420 20036 7472
rect 20904 7420 20956 7472
rect 21088 7420 21140 7472
rect 21640 7463 21692 7472
rect 21640 7429 21649 7463
rect 21649 7429 21683 7463
rect 21683 7429 21692 7463
rect 21640 7420 21692 7429
rect 16948 7352 17000 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17684 7352 17736 7404
rect 12992 7216 13044 7268
rect 14464 7284 14516 7336
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 13452 7148 13504 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14188 7259 14240 7268
rect 14188 7225 14197 7259
rect 14197 7225 14231 7259
rect 14231 7225 14240 7259
rect 14188 7216 14240 7225
rect 14556 7259 14608 7268
rect 14556 7225 14565 7259
rect 14565 7225 14599 7259
rect 14599 7225 14608 7259
rect 14556 7216 14608 7225
rect 18144 7352 18196 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 19248 7352 19300 7404
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 19524 7284 19576 7336
rect 20628 7352 20680 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 20904 7284 20956 7336
rect 16948 7216 17000 7268
rect 20168 7216 20220 7268
rect 15108 7148 15160 7200
rect 18880 7148 18932 7200
rect 20444 7148 20496 7200
rect 20996 7148 21048 7200
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 4169 7046 4221 7098
rect 4233 7046 4285 7098
rect 4297 7046 4349 7098
rect 4361 7046 4413 7098
rect 4425 7046 4477 7098
rect 10608 7046 10660 7098
rect 10672 7046 10724 7098
rect 10736 7046 10788 7098
rect 10800 7046 10852 7098
rect 10864 7046 10916 7098
rect 17047 7046 17099 7098
rect 17111 7046 17163 7098
rect 17175 7046 17227 7098
rect 17239 7046 17291 7098
rect 17303 7046 17355 7098
rect 23486 7046 23538 7098
rect 23550 7046 23602 7098
rect 23614 7046 23666 7098
rect 23678 7046 23730 7098
rect 23742 7046 23794 7098
rect 3240 6808 3292 6860
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 5448 6944 5500 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 8300 6944 8352 6996
rect 8760 6944 8812 6996
rect 9220 6944 9272 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 10416 6944 10468 6996
rect 11704 6944 11756 6996
rect 11980 6944 12032 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 20536 6987 20588 6996
rect 20536 6953 20545 6987
rect 20545 6953 20579 6987
rect 20579 6953 20588 6987
rect 20536 6944 20588 6953
rect 5448 6808 5500 6860
rect 3056 6672 3108 6724
rect 3700 6740 3752 6792
rect 3884 6740 3936 6792
rect 4804 6740 4856 6792
rect 5264 6740 5316 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 9128 6808 9180 6860
rect 9680 6808 9732 6860
rect 4160 6672 4212 6724
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4436 6715 4488 6724
rect 4436 6681 4445 6715
rect 4445 6681 4479 6715
rect 4479 6681 4488 6715
rect 4436 6672 4488 6681
rect 4712 6672 4764 6724
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10600 6876 10652 6928
rect 10968 6876 11020 6928
rect 11152 6876 11204 6928
rect 10232 6740 10284 6792
rect 10692 6740 10744 6792
rect 11796 6876 11848 6928
rect 13544 6876 13596 6928
rect 11612 6808 11664 6860
rect 20168 6876 20220 6928
rect 21456 6944 21508 6996
rect 11060 6672 11112 6724
rect 12440 6740 12492 6792
rect 16672 6808 16724 6860
rect 17408 6808 17460 6860
rect 13084 6740 13136 6792
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 16304 6740 16356 6792
rect 17684 6740 17736 6792
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 19984 6740 20036 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20996 6851 21048 6860
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 21456 6808 21508 6860
rect 5908 6604 5960 6656
rect 6000 6604 6052 6656
rect 8484 6604 8536 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12992 6672 13044 6724
rect 16948 6672 17000 6724
rect 17408 6672 17460 6724
rect 19156 6672 19208 6724
rect 21088 6740 21140 6792
rect 21916 6672 21968 6724
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 18052 6604 18104 6656
rect 19064 6604 19116 6656
rect 19984 6604 20036 6656
rect 4829 6502 4881 6554
rect 4893 6502 4945 6554
rect 4957 6502 5009 6554
rect 5021 6502 5073 6554
rect 5085 6502 5137 6554
rect 11268 6502 11320 6554
rect 11332 6502 11384 6554
rect 11396 6502 11448 6554
rect 11460 6502 11512 6554
rect 11524 6502 11576 6554
rect 17707 6502 17759 6554
rect 17771 6502 17823 6554
rect 17835 6502 17887 6554
rect 17899 6502 17951 6554
rect 17963 6502 18015 6554
rect 24146 6502 24198 6554
rect 24210 6502 24262 6554
rect 24274 6502 24326 6554
rect 24338 6502 24390 6554
rect 24402 6502 24454 6554
rect 940 6264 992 6316
rect 3884 6332 3936 6384
rect 4528 6400 4580 6452
rect 4804 6400 4856 6452
rect 5172 6400 5224 6452
rect 6092 6400 6144 6452
rect 9496 6400 9548 6452
rect 9956 6400 10008 6452
rect 10600 6400 10652 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 20076 6400 20128 6452
rect 21916 6443 21968 6452
rect 21916 6409 21925 6443
rect 21925 6409 21959 6443
rect 21959 6409 21968 6443
rect 21916 6400 21968 6409
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 5448 6332 5500 6384
rect 5908 6375 5960 6384
rect 5908 6341 5917 6375
rect 5917 6341 5951 6375
rect 5951 6341 5960 6375
rect 5908 6332 5960 6341
rect 3792 6196 3844 6248
rect 4436 6196 4488 6248
rect 5264 6264 5316 6316
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5724 6264 5776 6316
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 7288 6307 7340 6316
rect 6736 6264 6788 6273
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 8208 6332 8260 6384
rect 9128 6375 9180 6384
rect 9128 6341 9137 6375
rect 9137 6341 9171 6375
rect 9171 6341 9180 6375
rect 9128 6332 9180 6341
rect 9680 6332 9732 6384
rect 5724 6128 5776 6180
rect 6000 6128 6052 6180
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 6920 6196 6972 6248
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 6644 6060 6696 6112
rect 7472 6060 7524 6112
rect 8116 6060 8168 6112
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9220 6196 9272 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10140 6196 10192 6248
rect 10416 6196 10468 6248
rect 9772 6060 9824 6112
rect 10232 6060 10284 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 17408 6332 17460 6384
rect 18880 6332 18932 6384
rect 15384 6196 15436 6248
rect 18696 6264 18748 6316
rect 21088 6332 21140 6384
rect 18328 6196 18380 6248
rect 19984 6264 20036 6316
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 21456 6264 21508 6316
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 20720 6128 20772 6180
rect 20904 6171 20956 6180
rect 20904 6137 20913 6171
rect 20913 6137 20947 6171
rect 20947 6137 20956 6171
rect 20904 6128 20956 6137
rect 15016 6060 15068 6112
rect 19616 6060 19668 6112
rect 4169 5958 4221 6010
rect 4233 5958 4285 6010
rect 4297 5958 4349 6010
rect 4361 5958 4413 6010
rect 4425 5958 4477 6010
rect 10608 5958 10660 6010
rect 10672 5958 10724 6010
rect 10736 5958 10788 6010
rect 10800 5958 10852 6010
rect 10864 5958 10916 6010
rect 17047 5958 17099 6010
rect 17111 5958 17163 6010
rect 17175 5958 17227 6010
rect 17239 5958 17291 6010
rect 17303 5958 17355 6010
rect 23486 5958 23538 6010
rect 23550 5958 23602 6010
rect 23614 5958 23666 6010
rect 23678 5958 23730 6010
rect 23742 5958 23794 6010
rect 4620 5856 4672 5908
rect 5264 5856 5316 5908
rect 6276 5856 6328 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 10140 5856 10192 5908
rect 10324 5856 10376 5908
rect 12900 5856 12952 5908
rect 12992 5856 13044 5908
rect 6552 5788 6604 5840
rect 9864 5788 9916 5840
rect 5172 5720 5224 5772
rect 5356 5720 5408 5772
rect 5632 5695 5684 5704
rect 2228 5584 2280 5636
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 6920 5720 6972 5772
rect 13912 5788 13964 5840
rect 19340 5831 19392 5840
rect 19340 5797 19349 5831
rect 19349 5797 19383 5831
rect 19383 5797 19392 5831
rect 19340 5788 19392 5797
rect 5448 5584 5500 5636
rect 6000 5584 6052 5636
rect 6736 5652 6788 5704
rect 8944 5652 8996 5704
rect 9496 5652 9548 5704
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 16672 5652 16724 5704
rect 9220 5584 9272 5636
rect 7196 5516 7248 5568
rect 9496 5516 9548 5568
rect 9772 5584 9824 5636
rect 13360 5584 13412 5636
rect 15016 5584 15068 5636
rect 20076 5788 20128 5840
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20352 5720 20404 5772
rect 14372 5516 14424 5568
rect 19156 5584 19208 5636
rect 19432 5584 19484 5636
rect 18236 5516 18288 5568
rect 19524 5516 19576 5568
rect 26332 5652 26384 5704
rect 4829 5414 4881 5466
rect 4893 5414 4945 5466
rect 4957 5414 5009 5466
rect 5021 5414 5073 5466
rect 5085 5414 5137 5466
rect 11268 5414 11320 5466
rect 11332 5414 11384 5466
rect 11396 5414 11448 5466
rect 11460 5414 11512 5466
rect 11524 5414 11576 5466
rect 17707 5414 17759 5466
rect 17771 5414 17823 5466
rect 17835 5414 17887 5466
rect 17899 5414 17951 5466
rect 17963 5414 18015 5466
rect 24146 5414 24198 5466
rect 24210 5414 24262 5466
rect 24274 5414 24326 5466
rect 24338 5414 24390 5466
rect 24402 5414 24454 5466
rect 5632 5312 5684 5364
rect 6276 5312 6328 5364
rect 6920 5244 6972 5296
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 1584 5176 1636 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 9128 5176 9180 5228
rect 9496 5176 9548 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13084 5176 13136 5228
rect 13452 5176 13504 5228
rect 13636 5287 13688 5296
rect 13636 5253 13645 5287
rect 13645 5253 13679 5287
rect 13679 5253 13688 5287
rect 13636 5244 13688 5253
rect 9220 5108 9272 5160
rect 14004 5176 14056 5228
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 19340 5312 19392 5364
rect 16580 5176 16632 5228
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 19616 5176 19668 5228
rect 13912 5108 13964 5117
rect 12164 5040 12216 5092
rect 13268 5040 13320 5092
rect 18328 5108 18380 5160
rect 20904 5108 20956 5160
rect 21824 5108 21876 5160
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10508 4972 10560 5024
rect 13084 4972 13136 5024
rect 14004 4972 14056 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 15108 4972 15160 5024
rect 19248 4972 19300 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 4169 4870 4221 4922
rect 4233 4870 4285 4922
rect 4297 4870 4349 4922
rect 4361 4870 4413 4922
rect 4425 4870 4477 4922
rect 10608 4870 10660 4922
rect 10672 4870 10724 4922
rect 10736 4870 10788 4922
rect 10800 4870 10852 4922
rect 10864 4870 10916 4922
rect 17047 4870 17099 4922
rect 17111 4870 17163 4922
rect 17175 4870 17227 4922
rect 17239 4870 17291 4922
rect 17303 4870 17355 4922
rect 23486 4870 23538 4922
rect 23550 4870 23602 4922
rect 23614 4870 23666 4922
rect 23678 4870 23730 4922
rect 23742 4870 23794 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 10048 4768 10100 4820
rect 11060 4768 11112 4820
rect 6184 4632 6236 4684
rect 8300 4632 8352 4684
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 940 4564 992 4616
rect 4712 4564 4764 4616
rect 5172 4564 5224 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 8024 4564 8076 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 13084 4700 13136 4752
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 13544 4768 13596 4820
rect 15568 4768 15620 4820
rect 17408 4768 17460 4820
rect 20812 4768 20864 4820
rect 13912 4564 13964 4616
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 15108 4632 15160 4684
rect 16580 4632 16632 4684
rect 18236 4700 18288 4752
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15016 4564 15068 4616
rect 4436 4496 4488 4548
rect 5540 4539 5592 4548
rect 5540 4505 5549 4539
rect 5549 4505 5583 4539
rect 5583 4505 5592 4539
rect 5540 4496 5592 4505
rect 6276 4496 6328 4548
rect 4252 4428 4304 4480
rect 4528 4428 4580 4480
rect 9956 4471 10008 4480
rect 9956 4437 9965 4471
rect 9965 4437 9999 4471
rect 9999 4437 10008 4471
rect 9956 4428 10008 4437
rect 10232 4428 10284 4480
rect 12900 4496 12952 4548
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 12992 4428 13044 4480
rect 14372 4539 14424 4548
rect 14372 4505 14381 4539
rect 14381 4505 14415 4539
rect 14415 4505 14424 4539
rect 14372 4496 14424 4505
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 16764 4564 16816 4616
rect 17040 4675 17092 4684
rect 17040 4641 17049 4675
rect 17049 4641 17083 4675
rect 17083 4641 17092 4675
rect 17040 4632 17092 4641
rect 18052 4632 18104 4684
rect 19156 4632 19208 4684
rect 19432 4632 19484 4684
rect 18420 4564 18472 4616
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 18236 4539 18288 4548
rect 18236 4505 18245 4539
rect 18245 4505 18279 4539
rect 18279 4505 18288 4539
rect 18236 4496 18288 4505
rect 19984 4496 20036 4548
rect 13912 4428 13964 4437
rect 15660 4428 15712 4480
rect 16948 4428 17000 4480
rect 17224 4428 17276 4480
rect 18144 4428 18196 4480
rect 4829 4326 4881 4378
rect 4893 4326 4945 4378
rect 4957 4326 5009 4378
rect 5021 4326 5073 4378
rect 5085 4326 5137 4378
rect 11268 4326 11320 4378
rect 11332 4326 11384 4378
rect 11396 4326 11448 4378
rect 11460 4326 11512 4378
rect 11524 4326 11576 4378
rect 17707 4326 17759 4378
rect 17771 4326 17823 4378
rect 17835 4326 17887 4378
rect 17899 4326 17951 4378
rect 17963 4326 18015 4378
rect 24146 4326 24198 4378
rect 24210 4326 24262 4378
rect 24274 4326 24326 4378
rect 24338 4326 24390 4378
rect 24402 4326 24454 4378
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 10048 4224 10100 4276
rect 4160 4156 4212 4208
rect 3700 4088 3752 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 5172 4156 5224 4208
rect 6368 4156 6420 4208
rect 4712 4020 4764 4072
rect 5724 4131 5776 4140
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 8300 4156 8352 4208
rect 8852 4156 8904 4208
rect 12532 4224 12584 4276
rect 12624 4224 12676 4276
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 12992 4156 13044 4208
rect 4620 3952 4672 4004
rect 8024 4020 8076 4072
rect 8484 4020 8536 4072
rect 9772 4020 9824 4072
rect 11060 4020 11112 4072
rect 6644 3952 6696 4004
rect 9588 3952 9640 4004
rect 12440 4088 12492 4140
rect 12716 4088 12768 4140
rect 13360 4156 13412 4208
rect 13912 4224 13964 4276
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 14096 4156 14148 4208
rect 15476 4156 15528 4208
rect 13452 3952 13504 4004
rect 14924 4020 14976 4072
rect 3976 3884 4028 3936
rect 4160 3884 4212 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 6276 3884 6328 3936
rect 6736 3884 6788 3936
rect 9772 3884 9824 3936
rect 10416 3884 10468 3936
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 13360 3884 13412 3936
rect 14740 3884 14792 3936
rect 16212 4156 16264 4208
rect 16764 4199 16816 4208
rect 16764 4165 16773 4199
rect 16773 4165 16807 4199
rect 16807 4165 16816 4199
rect 16764 4156 16816 4165
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 18052 4224 18104 4276
rect 20444 4224 20496 4276
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 18144 4088 18196 4140
rect 18236 4088 18288 4140
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 16120 3952 16172 4004
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 17316 4020 17368 4072
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 16580 3952 16632 4004
rect 15476 3884 15528 3893
rect 17316 3884 17368 3936
rect 18420 3952 18472 4004
rect 19064 4088 19116 4140
rect 19248 4088 19300 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 26332 3995 26384 4004
rect 26332 3961 26341 3995
rect 26341 3961 26375 3995
rect 26375 3961 26384 3995
rect 26332 3952 26384 3961
rect 17684 3884 17736 3936
rect 4169 3782 4221 3834
rect 4233 3782 4285 3834
rect 4297 3782 4349 3834
rect 4361 3782 4413 3834
rect 4425 3782 4477 3834
rect 10608 3782 10660 3834
rect 10672 3782 10724 3834
rect 10736 3782 10788 3834
rect 10800 3782 10852 3834
rect 10864 3782 10916 3834
rect 17047 3782 17099 3834
rect 17111 3782 17163 3834
rect 17175 3782 17227 3834
rect 17239 3782 17291 3834
rect 17303 3782 17355 3834
rect 23486 3782 23538 3834
rect 23550 3782 23602 3834
rect 23614 3782 23666 3834
rect 23678 3782 23730 3834
rect 23742 3782 23794 3834
rect 5724 3680 5776 3732
rect 10232 3680 10284 3732
rect 12164 3680 12216 3732
rect 13544 3680 13596 3732
rect 16212 3680 16264 3732
rect 4068 3544 4120 3596
rect 6368 3544 6420 3596
rect 8300 3544 8352 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 12992 3544 13044 3596
rect 3700 3476 3752 3528
rect 4252 3476 4304 3528
rect 5724 3476 5776 3528
rect 8392 3476 8444 3528
rect 9588 3476 9640 3528
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 6920 3408 6972 3460
rect 8024 3408 8076 3460
rect 6368 3340 6420 3392
rect 7380 3340 7432 3392
rect 11612 3408 11664 3460
rect 12532 3408 12584 3460
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 16856 3544 16908 3596
rect 19064 3544 19116 3596
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 9128 3340 9180 3392
rect 13452 3451 13504 3460
rect 13452 3417 13461 3451
rect 13461 3417 13495 3451
rect 13495 3417 13504 3451
rect 13452 3408 13504 3417
rect 14372 3408 14424 3460
rect 14832 3408 14884 3460
rect 14096 3340 14148 3392
rect 18512 3383 18564 3392
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 4829 3238 4881 3290
rect 4893 3238 4945 3290
rect 4957 3238 5009 3290
rect 5021 3238 5073 3290
rect 5085 3238 5137 3290
rect 11268 3238 11320 3290
rect 11332 3238 11384 3290
rect 11396 3238 11448 3290
rect 11460 3238 11512 3290
rect 11524 3238 11576 3290
rect 17707 3238 17759 3290
rect 17771 3238 17823 3290
rect 17835 3238 17887 3290
rect 17899 3238 17951 3290
rect 17963 3238 18015 3290
rect 24146 3238 24198 3290
rect 24210 3238 24262 3290
rect 24274 3238 24326 3290
rect 24338 3238 24390 3290
rect 24402 3238 24454 3290
rect 6000 3136 6052 3188
rect 4068 3068 4120 3120
rect 4620 3068 4672 3120
rect 6184 3068 6236 3120
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8024 3136 8076 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 11060 3136 11112 3188
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 5816 2932 5868 2984
rect 6276 2932 6328 2984
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8392 3000 8444 3052
rect 9128 3068 9180 3120
rect 9772 3068 9824 3120
rect 8668 3000 8720 3052
rect 8944 3000 8996 3052
rect 15200 3000 15252 3052
rect 16856 3068 16908 3120
rect 16948 3111 17000 3120
rect 16948 3077 16957 3111
rect 16957 3077 16991 3111
rect 16991 3077 17000 3111
rect 16948 3068 17000 3077
rect 18512 3068 18564 3120
rect 5540 2864 5592 2916
rect 8300 2932 8352 2984
rect 9956 2932 10008 2984
rect 5724 2796 5776 2848
rect 6552 2796 6604 2848
rect 4169 2694 4221 2746
rect 4233 2694 4285 2746
rect 4297 2694 4349 2746
rect 4361 2694 4413 2746
rect 4425 2694 4477 2746
rect 10608 2694 10660 2746
rect 10672 2694 10724 2746
rect 10736 2694 10788 2746
rect 10800 2694 10852 2746
rect 10864 2694 10916 2746
rect 17047 2694 17099 2746
rect 17111 2694 17163 2746
rect 17175 2694 17227 2746
rect 17239 2694 17291 2746
rect 17303 2694 17355 2746
rect 23486 2694 23538 2746
rect 23550 2694 23602 2746
rect 23614 2694 23666 2746
rect 23678 2694 23730 2746
rect 23742 2694 23794 2746
rect 2412 2592 2464 2644
rect 5540 2592 5592 2644
rect 9772 2592 9824 2644
rect 940 2388 992 2440
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6644 2388 6696 2440
rect 10140 2456 10192 2508
rect 16304 2456 16356 2508
rect 8944 2388 8996 2440
rect 11152 2388 11204 2440
rect 14280 2388 14332 2440
rect 15844 2388 15896 2440
rect 6000 2320 6052 2372
rect 9956 2320 10008 2372
rect 13912 2320 13964 2372
rect 16396 2320 16448 2372
rect 18144 2295 18196 2304
rect 18144 2261 18153 2295
rect 18153 2261 18187 2295
rect 18187 2261 18196 2295
rect 18144 2252 18196 2261
rect 21824 2252 21876 2304
rect 25780 2252 25832 2304
rect 4829 2150 4881 2202
rect 4893 2150 4945 2202
rect 4957 2150 5009 2202
rect 5021 2150 5073 2202
rect 5085 2150 5137 2202
rect 11268 2150 11320 2202
rect 11332 2150 11384 2202
rect 11396 2150 11448 2202
rect 11460 2150 11512 2202
rect 11524 2150 11576 2202
rect 17707 2150 17759 2202
rect 17771 2150 17823 2202
rect 17835 2150 17887 2202
rect 17899 2150 17951 2202
rect 17963 2150 18015 2202
rect 24146 2150 24198 2202
rect 24210 2150 24262 2202
rect 24274 2150 24326 2202
rect 24338 2150 24390 2202
rect 24402 2150 24454 2202
<< metal2 >>
rect 3422 29332 3478 30132
rect 10414 29332 10470 30132
rect 17406 29332 17462 30132
rect 24398 29458 24454 30132
rect 24398 29430 24808 29458
rect 24398 29332 24454 29430
rect 2226 28112 2282 28121
rect 2226 28047 2282 28056
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24274 1440 24754
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 938 23760 994 23769
rect 938 23695 940 23704
rect 992 23695 994 23704
rect 940 23666 992 23672
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 938 21584 994 21593
rect 1412 21554 1440 24210
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 938 21519 994 21528
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21010 1440 21490
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1596 19961 1624 21830
rect 2240 20754 2268 28047
rect 3436 27606 3464 29332
rect 4169 27772 4477 27781
rect 4169 27770 4175 27772
rect 4231 27770 4255 27772
rect 4311 27770 4335 27772
rect 4391 27770 4415 27772
rect 4471 27770 4477 27772
rect 4231 27718 4233 27770
rect 4413 27718 4415 27770
rect 4169 27716 4175 27718
rect 4231 27716 4255 27718
rect 4311 27716 4335 27718
rect 4391 27716 4415 27718
rect 4471 27716 4477 27718
rect 4169 27707 4477 27716
rect 10428 27606 10456 29332
rect 10608 27772 10916 27781
rect 10608 27770 10614 27772
rect 10670 27770 10694 27772
rect 10750 27770 10774 27772
rect 10830 27770 10854 27772
rect 10910 27770 10916 27772
rect 10670 27718 10672 27770
rect 10852 27718 10854 27770
rect 10608 27716 10614 27718
rect 10670 27716 10694 27718
rect 10750 27716 10774 27718
rect 10830 27716 10854 27718
rect 10910 27716 10916 27718
rect 10608 27707 10916 27716
rect 17047 27772 17355 27781
rect 17047 27770 17053 27772
rect 17109 27770 17133 27772
rect 17189 27770 17213 27772
rect 17269 27770 17293 27772
rect 17349 27770 17355 27772
rect 17109 27718 17111 27770
rect 17291 27718 17293 27770
rect 17047 27716 17053 27718
rect 17109 27716 17133 27718
rect 17189 27716 17213 27718
rect 17269 27716 17293 27718
rect 17349 27716 17355 27718
rect 17047 27707 17355 27716
rect 17420 27606 17448 29332
rect 23486 27772 23794 27781
rect 23486 27770 23492 27772
rect 23548 27770 23572 27772
rect 23628 27770 23652 27772
rect 23708 27770 23732 27772
rect 23788 27770 23794 27772
rect 23548 27718 23550 27770
rect 23730 27718 23732 27770
rect 23486 27716 23492 27718
rect 23548 27716 23572 27718
rect 23628 27716 23652 27718
rect 23708 27716 23732 27718
rect 23788 27716 23794 27718
rect 23486 27707 23794 27716
rect 3424 27600 3476 27606
rect 3424 27542 3476 27548
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 24780 27554 24808 29430
rect 24860 27600 24912 27606
rect 24780 27548 24860 27554
rect 24780 27542 24912 27548
rect 24780 27526 24900 27542
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3344 26382 3372 26930
rect 3608 26784 3660 26790
rect 4172 26772 4200 27066
rect 4356 27062 4384 27270
rect 4829 27228 5137 27237
rect 4829 27226 4835 27228
rect 4891 27226 4915 27228
rect 4971 27226 4995 27228
rect 5051 27226 5075 27228
rect 5131 27226 5137 27228
rect 4891 27174 4893 27226
rect 5073 27174 5075 27226
rect 4829 27172 4835 27174
rect 4891 27172 4915 27174
rect 4971 27172 4995 27174
rect 5051 27172 5075 27174
rect 5131 27172 5137 27174
rect 4829 27163 5137 27172
rect 4344 27056 4396 27062
rect 4344 26998 4396 27004
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 3608 26726 3660 26732
rect 4080 26744 4200 26772
rect 3620 26382 3648 26726
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3804 26382 3832 26522
rect 3884 26512 3936 26518
rect 4080 26466 4108 26744
rect 4169 26684 4477 26693
rect 4169 26682 4175 26684
rect 4231 26682 4255 26684
rect 4311 26682 4335 26684
rect 4391 26682 4415 26684
rect 4471 26682 4477 26684
rect 4231 26630 4233 26682
rect 4413 26630 4415 26682
rect 4169 26628 4175 26630
rect 4231 26628 4255 26630
rect 4311 26628 4335 26630
rect 4391 26628 4415 26630
rect 4471 26628 4477 26630
rect 4169 26619 4477 26628
rect 3884 26454 3936 26460
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 3608 26376 3660 26382
rect 3608 26318 3660 26324
rect 3792 26376 3844 26382
rect 3792 26318 3844 26324
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3160 25906 3188 26182
rect 3422 25936 3478 25945
rect 3148 25900 3200 25906
rect 3422 25871 3478 25880
rect 3148 25842 3200 25848
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2976 24750 3004 25774
rect 3148 24880 3200 24886
rect 3148 24822 3200 24828
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 3160 24410 3188 24822
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 2792 23866 2820 24074
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2884 23730 2912 24142
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2792 23118 2820 23462
rect 2884 23186 2912 23666
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2884 22030 2912 23122
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2240 20726 2360 20754
rect 1582 19952 1638 19961
rect 1582 19887 1638 19896
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 1582 19816 1638 19825
rect 952 19417 980 19790
rect 1582 19751 1638 19760
rect 1596 19718 1624 19751
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 938 19408 994 19417
rect 938 19343 994 19352
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1504 18290 1532 18702
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 952 17241 980 17614
rect 938 17232 994 17241
rect 938 17167 994 17176
rect 1504 16658 1532 18226
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 17338 1624 17478
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1688 16114 1716 16594
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1596 15706 1624 15943
rect 2240 15706 2268 16458
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 12889 1440 13874
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13326 1716 13670
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1398 12880 1454 12889
rect 1872 12850 1900 13262
rect 1398 12815 1454 12824
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10713 1440 11086
rect 1872 10742 1900 12786
rect 2332 12238 2360 20726
rect 2424 19378 2452 21966
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2516 20874 2544 21830
rect 2792 21554 2820 21830
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2976 21010 3004 21830
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2792 18426 2820 19110
rect 2884 18766 2912 19450
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3160 18834 3188 19246
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3252 16402 3280 23054
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 3344 21690 3372 21966
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3344 19242 3372 19314
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 3344 18834 3372 19178
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3436 17882 3464 25871
rect 3896 25838 3924 26454
rect 3988 26438 4108 26466
rect 3988 26382 4016 26438
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 5172 26308 5224 26314
rect 5172 26250 5224 26256
rect 4829 26140 5137 26149
rect 4829 26138 4835 26140
rect 4891 26138 4915 26140
rect 4971 26138 4995 26140
rect 5051 26138 5075 26140
rect 5131 26138 5137 26140
rect 4891 26086 4893 26138
rect 5073 26086 5075 26138
rect 4829 26084 4835 26086
rect 4891 26084 4915 26086
rect 4971 26084 4995 26086
rect 5051 26084 5075 26086
rect 5131 26084 5137 26086
rect 4829 26075 5137 26084
rect 5184 26042 5212 26250
rect 5172 26036 5224 26042
rect 5172 25978 5224 25984
rect 3884 25832 3936 25838
rect 3884 25774 3936 25780
rect 5276 25702 5304 26862
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 4169 25596 4477 25605
rect 4169 25594 4175 25596
rect 4231 25594 4255 25596
rect 4311 25594 4335 25596
rect 4391 25594 4415 25596
rect 4471 25594 4477 25596
rect 4231 25542 4233 25594
rect 4413 25542 4415 25594
rect 4169 25540 4175 25542
rect 4231 25540 4255 25542
rect 4311 25540 4335 25542
rect 4391 25540 4415 25542
rect 4471 25540 4477 25542
rect 4169 25531 4477 25540
rect 4528 25492 4580 25498
rect 4528 25434 4580 25440
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 3608 25220 3660 25226
rect 3608 25162 3660 25168
rect 3620 24614 3648 25162
rect 4080 24818 4108 25298
rect 4540 25294 4568 25434
rect 5276 25294 5304 25638
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 4344 25152 4396 25158
rect 4344 25094 4396 25100
rect 4356 24886 4384 25094
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4344 24880 4396 24886
rect 4344 24822 4396 24828
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3620 24206 3648 24550
rect 3712 24274 3740 24550
rect 3896 24410 3924 24686
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 3988 23866 4016 24754
rect 4080 24342 4108 24754
rect 4344 24744 4396 24750
rect 4448 24732 4476 24890
rect 4396 24704 4476 24732
rect 4344 24686 4396 24692
rect 4169 24508 4477 24517
rect 4169 24506 4175 24508
rect 4231 24506 4255 24508
rect 4311 24506 4335 24508
rect 4391 24506 4415 24508
rect 4471 24506 4477 24508
rect 4231 24454 4233 24506
rect 4413 24454 4415 24506
rect 4169 24452 4175 24454
rect 4231 24452 4255 24454
rect 4311 24452 4335 24454
rect 4391 24452 4415 24454
rect 4471 24452 4477 24454
rect 4169 24443 4477 24452
rect 4068 24336 4120 24342
rect 4068 24278 4120 24284
rect 4540 24274 4568 25230
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4632 24886 4660 25094
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4528 24268 4580 24274
rect 4528 24210 4580 24216
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4172 23662 4200 24142
rect 4264 24070 4292 24142
rect 4632 24138 4660 24822
rect 4724 24818 4752 25162
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 4829 25052 5137 25061
rect 4829 25050 4835 25052
rect 4891 25050 4915 25052
rect 4971 25050 4995 25052
rect 5051 25050 5075 25052
rect 5131 25050 5137 25052
rect 4891 24998 4893 25050
rect 5073 24998 5075 25050
rect 4829 24996 4835 24998
rect 4891 24996 4915 24998
rect 4971 24996 4995 24998
rect 5051 24996 5075 24998
rect 5131 24996 5137 24998
rect 4829 24987 5137 24996
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4724 24188 4752 24754
rect 4816 24410 4844 24754
rect 5092 24750 5120 24822
rect 5184 24818 5212 25094
rect 5276 24818 5304 25230
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5080 24744 5132 24750
rect 5080 24686 5132 24692
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 4804 24200 4856 24206
rect 4724 24160 4804 24188
rect 4804 24142 4856 24148
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23798 4292 24006
rect 4252 23792 4304 23798
rect 4252 23734 4304 23740
rect 4632 23730 4660 24074
rect 4829 23964 5137 23973
rect 4829 23962 4835 23964
rect 4891 23962 4915 23964
rect 4971 23962 4995 23964
rect 5051 23962 5075 23964
rect 5131 23962 5137 23964
rect 4891 23910 4893 23962
rect 5073 23910 5075 23962
rect 4829 23908 4835 23910
rect 4891 23908 4915 23910
rect 4971 23908 4995 23910
rect 5051 23908 5075 23910
rect 5131 23908 5137 23910
rect 4829 23899 5137 23908
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4169 23420 4477 23429
rect 4169 23418 4175 23420
rect 4231 23418 4255 23420
rect 4311 23418 4335 23420
rect 4391 23418 4415 23420
rect 4471 23418 4477 23420
rect 4231 23366 4233 23418
rect 4413 23366 4415 23418
rect 4169 23364 4175 23366
rect 4231 23364 4255 23366
rect 4311 23364 4335 23366
rect 4391 23364 4415 23366
rect 4471 23364 4477 23366
rect 4169 23355 4477 23364
rect 4169 22332 4477 22341
rect 4169 22330 4175 22332
rect 4231 22330 4255 22332
rect 4311 22330 4335 22332
rect 4391 22330 4415 22332
rect 4471 22330 4477 22332
rect 4231 22278 4233 22330
rect 4413 22278 4415 22330
rect 4169 22276 4175 22278
rect 4231 22276 4255 22278
rect 4311 22276 4335 22278
rect 4391 22276 4415 22278
rect 4471 22276 4477 22278
rect 4169 22267 4477 22276
rect 4724 22234 4752 23598
rect 5276 23594 5304 24754
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 4829 22876 5137 22885
rect 4829 22874 4835 22876
rect 4891 22874 4915 22876
rect 4971 22874 4995 22876
rect 5051 22874 5075 22876
rect 5131 22874 5137 22876
rect 4891 22822 4893 22874
rect 5073 22822 5075 22874
rect 4829 22820 4835 22822
rect 4891 22820 4915 22822
rect 4971 22820 4995 22822
rect 5051 22820 5075 22822
rect 5131 22820 5137 22822
rect 4829 22811 5137 22820
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4068 22024 4120 22030
rect 4066 21992 4068 22001
rect 4160 22024 4212 22030
rect 4120 21992 4122 22001
rect 3516 21956 3568 21962
rect 4160 21966 4212 21972
rect 4066 21927 4122 21936
rect 3516 21898 3568 21904
rect 3528 21622 3556 21898
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3516 21616 3568 21622
rect 3568 21576 3648 21604
rect 3516 21558 3568 21564
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3528 20602 3556 21422
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3620 20330 3648 21576
rect 3712 20466 3740 21830
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3804 21350 3832 21626
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3804 20874 3832 21286
rect 3896 21146 3924 21422
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3804 20534 3832 20810
rect 3792 20528 3844 20534
rect 3792 20470 3844 20476
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 19378 3556 19654
rect 3896 19446 3924 21082
rect 3988 20602 4016 21490
rect 4172 21434 4200 21966
rect 4356 21486 4384 22170
rect 5368 22094 5396 27338
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 5448 26852 5500 26858
rect 5448 26794 5500 26800
rect 5460 26586 5488 26794
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5460 25430 5488 26522
rect 6000 25900 6052 25906
rect 6000 25842 6052 25848
rect 6012 25430 6040 25842
rect 5448 25424 5500 25430
rect 5448 25366 5500 25372
rect 6000 25424 6052 25430
rect 6000 25366 6052 25372
rect 5460 24206 5488 25366
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5552 24410 5580 24686
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5552 23866 5580 24346
rect 5644 24070 5672 24686
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 6012 23050 6040 25366
rect 6380 24818 6408 26930
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 25974 6500 26318
rect 6460 25968 6512 25974
rect 6460 25910 6512 25916
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6196 24342 6224 24754
rect 6564 24410 6592 24754
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6184 24336 6236 24342
rect 6184 24278 6236 24284
rect 6656 23730 6684 26386
rect 6748 24954 6776 26862
rect 6932 25702 6960 26930
rect 7024 25770 7052 27338
rect 7116 26466 7144 27338
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 7208 26586 7236 26930
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 7116 26438 7236 26466
rect 7208 26382 7236 26438
rect 7300 26382 7328 26726
rect 8116 26512 8168 26518
rect 8116 26454 8168 26460
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7208 26042 7236 26318
rect 7380 26240 7432 26246
rect 7380 26182 7432 26188
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 7012 25764 7064 25770
rect 7012 25706 7064 25712
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 7116 25498 7144 25910
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6748 23730 6776 24550
rect 6840 24070 6868 25094
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7024 24410 7052 24686
rect 7116 24614 7144 25434
rect 7208 25226 7236 25978
rect 7392 25974 7420 26182
rect 7380 25968 7432 25974
rect 7380 25910 7432 25916
rect 7392 25838 7420 25910
rect 7564 25900 7616 25906
rect 7616 25860 7696 25888
rect 7564 25842 7616 25848
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7392 25344 7420 25774
rect 7392 25316 7512 25344
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7392 24818 7420 25162
rect 7484 24818 7512 25316
rect 7668 25294 7696 25860
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7668 24818 7696 25230
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7116 24206 7144 24550
rect 7392 24206 7420 24754
rect 7668 24410 7696 24754
rect 8128 24750 8156 26454
rect 9140 26382 9168 26930
rect 10324 26784 10376 26790
rect 10324 26726 10376 26732
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9140 25430 9168 26318
rect 10336 26314 10364 26726
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9692 25498 9720 25910
rect 10232 25832 10284 25838
rect 10232 25774 10284 25780
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9128 25424 9180 25430
rect 9128 25366 9180 25372
rect 10244 25158 10272 25774
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7760 24274 7788 24550
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6182 23216 6238 23225
rect 6182 23151 6238 23160
rect 6196 23118 6224 23151
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6000 23044 6052 23050
rect 6000 22986 6052 22992
rect 6288 22098 6316 23666
rect 7116 23322 7144 23734
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 5184 22066 5396 22094
rect 6276 22092 6328 22098
rect 5080 22024 5132 22030
rect 5078 21992 5080 22001
rect 5132 21992 5134 22001
rect 4448 21950 4660 21978
rect 4448 21894 4476 21950
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4080 21406 4200 21434
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4080 21026 4108 21406
rect 4356 21350 4384 21422
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4169 21244 4477 21253
rect 4169 21242 4175 21244
rect 4231 21242 4255 21244
rect 4311 21242 4335 21244
rect 4391 21242 4415 21244
rect 4471 21242 4477 21244
rect 4231 21190 4233 21242
rect 4413 21190 4415 21242
rect 4169 21188 4175 21190
rect 4231 21188 4255 21190
rect 4311 21188 4335 21190
rect 4391 21188 4415 21190
rect 4471 21188 4477 21190
rect 4169 21179 4477 21188
rect 4160 21072 4212 21078
rect 4080 21020 4160 21026
rect 4080 21014 4212 21020
rect 4080 20998 4200 21014
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 4172 20398 4200 20998
rect 4632 20874 4660 21950
rect 5078 21927 5134 21936
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21622 4752 21830
rect 4829 21788 5137 21797
rect 4829 21786 4835 21788
rect 4891 21786 4915 21788
rect 4971 21786 4995 21788
rect 5051 21786 5075 21788
rect 5131 21786 5137 21788
rect 4891 21734 4893 21786
rect 5073 21734 5075 21786
rect 4829 21732 4835 21734
rect 4891 21732 4915 21734
rect 4971 21732 4995 21734
rect 5051 21732 5075 21734
rect 5131 21732 5137 21734
rect 4829 21723 5137 21732
rect 4712 21616 4764 21622
rect 5184 21604 5212 22066
rect 6276 22034 6328 22040
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5908 22024 5960 22030
rect 6288 22003 6316 22034
rect 5908 21966 5960 21972
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5092 21576 5212 21604
rect 4764 21564 4844 21570
rect 4712 21558 4844 21564
rect 4724 21542 4844 21558
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4724 20602 4752 21422
rect 4816 20942 4844 21542
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4908 21146 4936 21286
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 5092 20856 5120 21576
rect 5172 21538 5224 21544
rect 5172 21480 5224 21486
rect 5184 21146 5212 21480
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5276 21078 5304 21830
rect 5368 21554 5396 21830
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5460 21434 5488 21898
rect 5368 21406 5488 21434
rect 5368 21350 5396 21406
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5368 21146 5396 21286
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5092 20828 5304 20856
rect 4829 20700 5137 20709
rect 4829 20698 4835 20700
rect 4891 20698 4915 20700
rect 4971 20698 4995 20700
rect 5051 20698 5075 20700
rect 5131 20698 5137 20700
rect 4891 20646 4893 20698
rect 5073 20646 5075 20698
rect 4829 20644 4835 20646
rect 4891 20644 4915 20646
rect 4971 20644 4995 20646
rect 5051 20644 5075 20646
rect 5131 20644 5137 20646
rect 4829 20635 5137 20644
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 4080 19242 4108 20266
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4169 20156 4477 20165
rect 4169 20154 4175 20156
rect 4231 20154 4255 20156
rect 4311 20154 4335 20156
rect 4391 20154 4415 20156
rect 4471 20154 4477 20156
rect 4231 20102 4233 20154
rect 4413 20102 4415 20154
rect 4169 20100 4175 20102
rect 4231 20100 4255 20102
rect 4311 20100 4335 20102
rect 4391 20100 4415 20102
rect 4471 20100 4477 20102
rect 4169 20091 4477 20100
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4172 19378 4200 19450
rect 4540 19378 4568 20198
rect 5184 19854 5212 20470
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4169 19068 4477 19077
rect 4169 19066 4175 19068
rect 4231 19066 4255 19068
rect 4311 19066 4335 19068
rect 4391 19066 4415 19068
rect 4471 19066 4477 19068
rect 4231 19014 4233 19066
rect 4413 19014 4415 19066
rect 4169 19012 4175 19014
rect 4231 19012 4255 19014
rect 4311 19012 4335 19014
rect 4391 19012 4415 19014
rect 4471 19012 4477 19014
rect 4169 19003 4477 19012
rect 4540 18766 4568 19314
rect 4632 18834 4660 19790
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4724 19394 4752 19722
rect 4829 19612 5137 19621
rect 4829 19610 4835 19612
rect 4891 19610 4915 19612
rect 4971 19610 4995 19612
rect 5051 19610 5075 19612
rect 5131 19610 5137 19612
rect 4891 19558 4893 19610
rect 5073 19558 5075 19610
rect 4829 19556 4835 19558
rect 4891 19556 4915 19558
rect 4971 19556 4995 19558
rect 5051 19556 5075 19558
rect 5131 19556 5137 19558
rect 4829 19547 5137 19556
rect 5276 19417 5304 20828
rect 5368 19514 5396 20878
rect 5552 20602 5580 21966
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5644 21010 5672 21286
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5632 20528 5684 20534
rect 5632 20470 5684 20476
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5460 19854 5488 20266
rect 5644 20262 5672 20470
rect 5736 20466 5764 21490
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5828 20262 5856 21286
rect 5920 20806 5948 21966
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6196 21690 6224 21898
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21690 6500 21830
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6564 21570 6592 22714
rect 6472 21542 6592 21570
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 6012 20466 6040 21422
rect 6472 21418 6500 21542
rect 6552 21480 6604 21486
rect 6748 21434 6776 23122
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 21554 6868 21830
rect 7116 21554 7144 23054
rect 8036 23050 8064 24686
rect 8128 23254 8156 24686
rect 8220 24206 8248 24686
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8220 23866 8248 24142
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 8220 22710 8248 23802
rect 9312 23792 9364 23798
rect 9310 23760 9312 23769
rect 9364 23760 9366 23769
rect 9220 23724 9272 23730
rect 9310 23695 9366 23704
rect 9220 23666 9272 23672
rect 9034 23352 9090 23361
rect 9034 23287 9090 23296
rect 9128 23316 9180 23322
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8392 23112 8444 23118
rect 8956 23089 8984 23190
rect 9048 23186 9076 23287
rect 9128 23258 9180 23264
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 8392 23054 8444 23060
rect 8942 23080 8998 23089
rect 8208 22704 8260 22710
rect 8208 22646 8260 22652
rect 8404 22642 8432 23054
rect 8942 23015 8998 23024
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 8864 22642 8892 22918
rect 9140 22681 9168 23258
rect 9126 22672 9182 22681
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8852 22636 8904 22642
rect 9126 22607 9182 22616
rect 8852 22578 8904 22584
rect 8404 22030 8432 22578
rect 9140 22438 9168 22607
rect 9232 22574 9260 23666
rect 9968 23662 9996 24006
rect 10244 23866 10272 25094
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10322 23760 10378 23769
rect 10322 23695 10324 23704
rect 10376 23695 10378 23704
rect 10324 23666 10376 23672
rect 9772 23656 9824 23662
rect 9770 23624 9772 23633
rect 9956 23656 10008 23662
rect 9824 23624 9826 23633
rect 9956 23598 10008 23604
rect 9770 23559 9826 23568
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9220 22568 9272 22574
rect 9272 22528 9352 22556
rect 9220 22510 9272 22516
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22234 9168 22374
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9140 22098 9168 22170
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7208 21690 7236 21898
rect 9324 21876 9352 22528
rect 9416 22030 9444 23258
rect 9588 23180 9640 23186
rect 9508 23140 9588 23168
rect 9508 22574 9536 23140
rect 9588 23122 9640 23128
rect 9692 22760 9720 23462
rect 9862 23352 9918 23361
rect 9862 23287 9918 23296
rect 9876 23186 9904 23287
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9772 23112 9824 23118
rect 9770 23080 9772 23089
rect 9824 23080 9826 23089
rect 9770 23015 9826 23024
rect 9600 22732 9720 22760
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9508 22166 9536 22510
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9324 21848 9444 21876
rect 9416 21842 9444 21848
rect 9508 21842 9536 21898
rect 9416 21814 9536 21842
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6604 21428 6868 21434
rect 6552 21422 6868 21428
rect 6460 21412 6512 21418
rect 6564 21406 6868 21422
rect 6460 21354 6512 21360
rect 6840 21350 6868 21406
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6472 20466 6500 20742
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5828 19854 5856 20198
rect 6748 20058 6776 20334
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6840 19938 6868 21286
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6748 19910 6868 19938
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5262 19408 5318 19417
rect 4724 19366 4844 19394
rect 4816 19310 4844 19366
rect 5262 19343 5318 19352
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4816 18834 4844 19246
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 5460 18766 5488 19790
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 18358 3924 18566
rect 4829 18524 5137 18533
rect 4829 18522 4835 18524
rect 4891 18522 4915 18524
rect 4971 18522 4995 18524
rect 5051 18522 5075 18524
rect 5131 18522 5137 18524
rect 4891 18470 4893 18522
rect 5073 18470 5075 18522
rect 4829 18468 4835 18470
rect 4891 18468 4915 18470
rect 4971 18468 4995 18470
rect 5051 18468 5075 18470
rect 5131 18468 5137 18470
rect 4829 18459 5137 18468
rect 5184 18426 5212 18702
rect 5552 18698 5580 19790
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 5736 18970 5764 19314
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 3884 18352 3936 18358
rect 3884 18294 3936 18300
rect 4169 17980 4477 17989
rect 4169 17978 4175 17980
rect 4231 17978 4255 17980
rect 4311 17978 4335 17980
rect 4391 17978 4415 17980
rect 4471 17978 4477 17980
rect 4231 17926 4233 17978
rect 4413 17926 4415 17978
rect 4169 17924 4175 17926
rect 4231 17924 4255 17926
rect 4311 17924 4335 17926
rect 4391 17924 4415 17926
rect 4471 17924 4477 17926
rect 4169 17915 4477 17924
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 6288 17542 6316 19314
rect 6748 19310 6776 19910
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6932 18970 6960 19382
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 4829 17436 5137 17445
rect 4829 17434 4835 17436
rect 4891 17434 4915 17436
rect 4971 17434 4995 17436
rect 5051 17434 5075 17436
rect 5131 17434 5137 17436
rect 4891 17382 4893 17434
rect 5073 17382 5075 17434
rect 4829 17380 4835 17382
rect 4891 17380 4915 17382
rect 4971 17380 4995 17382
rect 5051 17380 5075 17382
rect 5131 17380 5137 17382
rect 4829 17371 5137 17380
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 2884 15638 2912 16390
rect 3160 15706 3188 16390
rect 3252 16374 3556 16402
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 15162 2820 15302
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2884 14822 2912 15574
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3344 15366 3372 15506
rect 3436 15502 3464 15846
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 3068 14482 3096 15030
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13734 2820 14214
rect 3160 14006 3188 15098
rect 3344 14550 3372 15302
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3436 14482 3464 15438
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 3252 13530 3280 14350
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3252 13326 3280 13466
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 2700 12374 2728 13262
rect 3344 12850 3372 14214
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 12986 3464 13806
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 3436 12306 3464 12786
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 1860 10736 1912 10742
rect 1398 10704 1454 10713
rect 1860 10678 1912 10684
rect 1398 10639 1454 10648
rect 1872 10130 1900 10678
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 9586 1900 10066
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 952 8537 980 8910
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 938 6352 994 6361
rect 938 6287 940 6296
rect 992 6287 994 6296
rect 940 6258 992 6264
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4826 1624 5170
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 952 2009 980 2382
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 2056 800 2084 12174
rect 3528 11286 3556 16374
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 15706 3648 15846
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3804 15094 3832 16458
rect 3896 15706 3924 17138
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16590 4108 16934
rect 4169 16892 4477 16901
rect 4169 16890 4175 16892
rect 4231 16890 4255 16892
rect 4311 16890 4335 16892
rect 4391 16890 4415 16892
rect 4471 16890 4477 16892
rect 4231 16838 4233 16890
rect 4413 16838 4415 16890
rect 4169 16836 4175 16838
rect 4231 16836 4255 16838
rect 4311 16836 4335 16838
rect 4391 16836 4415 16838
rect 4471 16836 4477 16838
rect 4169 16827 4477 16836
rect 4816 16794 4844 17138
rect 5092 16794 5120 17138
rect 6288 17134 6316 17478
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16794 5580 16934
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 6288 16658 6316 17070
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 5092 16454 5120 16526
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4829 16348 5137 16357
rect 4829 16346 4835 16348
rect 4891 16346 4915 16348
rect 4971 16346 4995 16348
rect 5051 16346 5075 16348
rect 5131 16346 5137 16348
rect 4891 16294 4893 16346
rect 5073 16294 5075 16346
rect 4829 16292 4835 16294
rect 4891 16292 4915 16294
rect 4971 16292 4995 16294
rect 5051 16292 5075 16294
rect 5131 16292 5137 16294
rect 4829 16283 5137 16292
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3712 14074 3740 14486
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3804 13138 3832 15030
rect 3896 14822 3924 15506
rect 3988 15162 4016 16118
rect 5184 16114 5212 16390
rect 6288 16182 6316 16594
rect 6656 16522 6684 17818
rect 7024 17678 7052 20810
rect 7116 19854 7144 21490
rect 8220 20602 8248 21626
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7300 20058 7328 20470
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 8404 19922 8432 20198
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8680 19854 8708 20742
rect 8956 20602 8984 20946
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 7116 18902 7144 19790
rect 8956 19786 8984 20538
rect 9048 19854 9076 20810
rect 9416 20058 9444 20946
rect 9600 20058 9628 22732
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9692 22545 9720 22578
rect 9772 22568 9824 22574
rect 9678 22536 9734 22545
rect 9772 22510 9824 22516
rect 9678 22471 9734 22480
rect 9680 21888 9732 21894
rect 9784 21876 9812 22510
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 22234 9904 22442
rect 9968 22234 9996 23598
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9956 22024 10008 22030
rect 9862 21992 9918 22001
rect 9956 21966 10008 21972
rect 9862 21927 9864 21936
rect 9916 21927 9918 21936
rect 9864 21898 9916 21904
rect 9732 21848 9812 21876
rect 9680 21830 9732 21836
rect 9968 21146 9996 21966
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9692 20466 9720 20878
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9784 20602 9812 20742
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8772 19378 8800 19654
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 8772 18766 8800 19314
rect 9048 18970 9076 19790
rect 9416 19514 9444 19994
rect 9876 19990 9904 20742
rect 9968 20466 9996 20810
rect 10060 20602 10088 22374
rect 10152 21894 10180 22578
rect 10244 22094 10272 22918
rect 10428 22522 10456 27338
rect 11268 27228 11576 27237
rect 11268 27226 11274 27228
rect 11330 27226 11354 27228
rect 11410 27226 11434 27228
rect 11490 27226 11514 27228
rect 11570 27226 11576 27228
rect 11330 27174 11332 27226
rect 11512 27174 11514 27226
rect 11268 27172 11274 27174
rect 11330 27172 11354 27174
rect 11410 27172 11434 27174
rect 11490 27172 11514 27174
rect 11570 27172 11576 27174
rect 11268 27163 11576 27172
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 10608 26684 10916 26693
rect 10608 26682 10614 26684
rect 10670 26682 10694 26684
rect 10750 26682 10774 26684
rect 10830 26682 10854 26684
rect 10910 26682 10916 26684
rect 10670 26630 10672 26682
rect 10852 26630 10854 26682
rect 10608 26628 10614 26630
rect 10670 26628 10694 26630
rect 10750 26628 10774 26630
rect 10830 26628 10854 26630
rect 10910 26628 10916 26630
rect 10608 26619 10916 26628
rect 10888 26438 11100 26466
rect 10888 26382 10916 26438
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 10796 25906 10824 26182
rect 10980 25974 11008 26318
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10608 25596 10916 25605
rect 10608 25594 10614 25596
rect 10670 25594 10694 25596
rect 10750 25594 10774 25596
rect 10830 25594 10854 25596
rect 10910 25594 10916 25596
rect 10670 25542 10672 25594
rect 10852 25542 10854 25594
rect 10608 25540 10614 25542
rect 10670 25540 10694 25542
rect 10750 25540 10774 25542
rect 10830 25540 10854 25542
rect 10910 25540 10916 25542
rect 10608 25531 10916 25540
rect 10980 25294 11008 25774
rect 11072 25702 11100 26438
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11268 26140 11576 26149
rect 11268 26138 11274 26140
rect 11330 26138 11354 26140
rect 11410 26138 11434 26140
rect 11490 26138 11514 26140
rect 11570 26138 11576 26140
rect 11330 26086 11332 26138
rect 11512 26086 11514 26138
rect 11268 26084 11274 26086
rect 11330 26084 11354 26086
rect 11410 26084 11434 26086
rect 11490 26084 11514 26086
rect 11570 26084 11576 26086
rect 11268 26075 11576 26084
rect 11624 26042 11652 26250
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 11716 25838 11744 25978
rect 11992 25974 12020 26930
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 12084 26314 12112 26726
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 12268 26042 12296 26862
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 11980 25968 12032 25974
rect 11900 25928 11980 25956
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11520 25764 11572 25770
rect 11520 25706 11572 25712
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11532 25498 11560 25706
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11268 25052 11576 25061
rect 11268 25050 11274 25052
rect 11330 25050 11354 25052
rect 11410 25050 11434 25052
rect 11490 25050 11514 25052
rect 11570 25050 11576 25052
rect 11330 24998 11332 25050
rect 11512 24998 11514 25050
rect 11268 24996 11274 24998
rect 11330 24996 11354 24998
rect 11410 24996 11434 24998
rect 11490 24996 11514 24998
rect 11570 24996 11576 24998
rect 11268 24987 11576 24996
rect 11716 24886 11744 25230
rect 11808 24954 11836 25842
rect 11900 25226 11928 25928
rect 11980 25910 12032 25916
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 12072 25832 12124 25838
rect 12072 25774 12124 25780
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11992 24954 12020 25774
rect 12084 25498 12112 25774
rect 12176 25498 12204 25910
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11704 24880 11756 24886
rect 11704 24822 11756 24828
rect 10608 24508 10916 24517
rect 10608 24506 10614 24508
rect 10670 24506 10694 24508
rect 10750 24506 10774 24508
rect 10830 24506 10854 24508
rect 10910 24506 10916 24508
rect 10670 24454 10672 24506
rect 10852 24454 10854 24506
rect 10608 24452 10614 24454
rect 10670 24452 10694 24454
rect 10750 24452 10774 24454
rect 10830 24452 10854 24454
rect 10910 24452 10916 24454
rect 10608 24443 10916 24452
rect 11060 24336 11112 24342
rect 11060 24278 11112 24284
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10520 23322 10548 23802
rect 10600 23656 10652 23662
rect 10598 23624 10600 23633
rect 10652 23624 10654 23633
rect 10704 23594 10732 24074
rect 10598 23559 10654 23568
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10608 23420 10916 23429
rect 10608 23418 10614 23420
rect 10670 23418 10694 23420
rect 10750 23418 10774 23420
rect 10830 23418 10854 23420
rect 10910 23418 10916 23420
rect 10670 23366 10672 23418
rect 10852 23366 10854 23418
rect 10608 23364 10614 23366
rect 10670 23364 10694 23366
rect 10750 23364 10774 23366
rect 10830 23364 10854 23366
rect 10910 23364 10916 23366
rect 10608 23355 10916 23364
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10336 22494 10456 22522
rect 10336 22234 10364 22494
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10244 22066 10364 22094
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10244 21690 10272 21898
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10336 21078 10364 22066
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9508 19378 9536 19722
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19378 9628 19654
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9232 18766 9260 19314
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9404 18760 9456 18766
rect 9508 18748 9536 19314
rect 9600 18766 9628 19314
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9456 18720 9536 18748
rect 9588 18760 9640 18766
rect 9404 18702 9456 18708
rect 9588 18702 9640 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 8312 17202 8340 18566
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9416 17338 9444 17614
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16794 8340 17138
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6564 16250 6592 16458
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4080 15570 4108 15914
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4169 15804 4477 15813
rect 4169 15802 4175 15804
rect 4231 15802 4255 15804
rect 4311 15802 4335 15804
rect 4391 15802 4415 15804
rect 4471 15802 4477 15804
rect 4231 15750 4233 15802
rect 4413 15750 4415 15802
rect 4169 15748 4175 15750
rect 4231 15748 4255 15750
rect 4311 15748 4335 15750
rect 4391 15748 4415 15750
rect 4471 15748 4477 15750
rect 4169 15739 4477 15748
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4356 15450 4384 15506
rect 4540 15502 4568 15846
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4080 15422 4384 15450
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 13258 3924 14758
rect 3988 14414 4016 15098
rect 4080 15094 4108 15422
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4169 14716 4477 14725
rect 4169 14714 4175 14716
rect 4231 14714 4255 14716
rect 4311 14714 4335 14716
rect 4391 14714 4415 14716
rect 4471 14714 4477 14716
rect 4231 14662 4233 14714
rect 4413 14662 4415 14714
rect 4169 14660 4175 14662
rect 4231 14660 4255 14662
rect 4311 14660 4335 14662
rect 4391 14660 4415 14662
rect 4471 14660 4477 14662
rect 4169 14651 4477 14660
rect 4632 14414 4660 15574
rect 4829 15260 5137 15269
rect 4829 15258 4835 15260
rect 4891 15258 4915 15260
rect 4971 15258 4995 15260
rect 5051 15258 5075 15260
rect 5131 15258 5137 15260
rect 4891 15206 4893 15258
rect 5073 15206 5075 15258
rect 4829 15204 4835 15206
rect 4891 15204 4915 15206
rect 4971 15204 4995 15206
rect 5051 15204 5075 15206
rect 5131 15204 5137 15206
rect 4829 15195 5137 15204
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3988 13802 4016 14214
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13818 4108 13874
rect 4172 13818 4200 14350
rect 4264 14074 4292 14350
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 4080 13790 4200 13818
rect 4724 13818 4752 14214
rect 4829 14172 5137 14181
rect 4829 14170 4835 14172
rect 4891 14170 4915 14172
rect 4971 14170 4995 14172
rect 5051 14170 5075 14172
rect 5131 14170 5137 14172
rect 4891 14118 4893 14170
rect 5073 14118 5075 14170
rect 4829 14116 4835 14118
rect 4891 14116 4915 14118
rect 4971 14116 4995 14118
rect 5051 14116 5075 14118
rect 5131 14116 5137 14118
rect 4829 14107 5137 14116
rect 5184 13938 5212 16050
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15434 5672 15846
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5736 15162 5764 16050
rect 6288 15502 6316 16118
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 15570 6592 16050
rect 6932 15978 6960 16186
rect 7300 16182 7328 16390
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 7208 15586 7236 16118
rect 7300 15978 7328 16118
rect 7392 16017 7420 16118
rect 7760 16046 7788 16390
rect 8404 16250 8432 16934
rect 8496 16794 8524 17070
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8588 16726 8616 17002
rect 9232 16794 9260 17070
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 7748 16040 7800 16046
rect 7378 16008 7434 16017
rect 7288 15972 7340 15978
rect 7748 15982 7800 15988
rect 7378 15943 7434 15952
rect 7288 15914 7340 15920
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 6552 15564 6604 15570
rect 7208 15558 7328 15586
rect 6552 15506 6604 15512
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4528 13796 4580 13802
rect 3988 13530 4016 13738
rect 3976 13524 4028 13530
rect 4080 13512 4108 13790
rect 4724 13790 4936 13818
rect 4528 13738 4580 13744
rect 4169 13628 4477 13637
rect 4169 13626 4175 13628
rect 4231 13626 4255 13628
rect 4311 13626 4335 13628
rect 4391 13626 4415 13628
rect 4471 13626 4477 13628
rect 4231 13574 4233 13626
rect 4413 13574 4415 13626
rect 4169 13572 4175 13574
rect 4231 13572 4255 13574
rect 4311 13572 4335 13574
rect 4391 13572 4415 13574
rect 4471 13572 4477 13574
rect 4169 13563 4477 13572
rect 4160 13524 4212 13530
rect 4080 13484 4160 13512
rect 3976 13466 4028 13472
rect 4160 13466 4212 13472
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3804 13110 3924 13138
rect 3896 12986 3924 13110
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3804 12238 3832 12922
rect 3976 12912 4028 12918
rect 3974 12880 3976 12889
rect 4028 12880 4030 12889
rect 3974 12815 4030 12824
rect 4172 12730 4200 13330
rect 4356 12918 4384 13398
rect 4540 13376 4568 13738
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4448 13348 4568 13376
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4080 12702 4200 12730
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12442 4016 12582
rect 3976 12436 4028 12442
rect 4080 12434 4108 12702
rect 4448 12646 4476 13348
rect 4632 12850 4660 13670
rect 4724 12850 4752 13670
rect 4908 13326 4936 13790
rect 5000 13530 5028 13874
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4896 13320 4948 13326
rect 5080 13320 5132 13326
rect 4896 13262 4948 13268
rect 5078 13288 5080 13297
rect 5132 13288 5134 13297
rect 5078 13223 5134 13232
rect 4829 13084 5137 13093
rect 4829 13082 4835 13084
rect 4891 13082 4915 13084
rect 4971 13082 4995 13084
rect 5051 13082 5075 13084
rect 5131 13082 5137 13084
rect 4891 13030 4893 13082
rect 5073 13030 5075 13082
rect 4829 13028 4835 13030
rect 4891 13028 4915 13030
rect 4971 13028 4995 13030
rect 5051 13028 5075 13030
rect 5131 13028 5137 13030
rect 4829 13019 5137 13028
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4169 12540 4477 12549
rect 4169 12538 4175 12540
rect 4231 12538 4255 12540
rect 4311 12538 4335 12540
rect 4391 12538 4415 12540
rect 4471 12538 4477 12540
rect 4231 12486 4233 12538
rect 4413 12486 4415 12538
rect 4169 12484 4175 12486
rect 4231 12484 4255 12486
rect 4311 12484 4335 12486
rect 4391 12484 4415 12486
rect 4471 12484 4477 12486
rect 4169 12475 4477 12484
rect 4540 12442 4568 12786
rect 5184 12714 5212 13670
rect 5276 13326 5304 14282
rect 6564 14074 6592 15506
rect 7300 15502 7328 15558
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15026 6684 15302
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 7300 14958 7328 15438
rect 7392 15366 7420 15846
rect 7668 15502 7696 15846
rect 7760 15502 7788 15846
rect 8496 15706 8524 16594
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8588 15706 8616 16050
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6656 13938 6684 14214
rect 6932 14074 6960 14894
rect 7392 14414 7420 15302
rect 7760 14414 7788 15302
rect 8496 14482 8524 15438
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 7208 14074 7236 14350
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 7116 13870 7144 13942
rect 7484 13938 7512 14214
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12918 5304 13262
rect 5460 13258 5488 13670
rect 5552 13530 5580 13806
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5460 12850 5488 13194
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5644 12782 5672 13330
rect 6472 13326 6500 13670
rect 7116 13530 7144 13806
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 4632 12442 4660 12650
rect 4528 12436 4580 12442
rect 4080 12406 4200 12434
rect 3976 12378 4028 12384
rect 4172 12306 4200 12406
rect 4528 12378 4580 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 5828 12374 5856 13262
rect 7116 12850 7144 13466
rect 7484 13326 7512 13874
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7576 13530 7604 13738
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 4829 11996 5137 12005
rect 4829 11994 4835 11996
rect 4891 11994 4915 11996
rect 4971 11994 4995 11996
rect 5051 11994 5075 11996
rect 5131 11994 5137 11996
rect 4891 11942 4893 11994
rect 5073 11942 5075 11994
rect 4829 11940 4835 11942
rect 4891 11940 4915 11942
rect 4971 11940 4995 11942
rect 5051 11940 5075 11942
rect 5131 11940 5137 11942
rect 4829 11931 5137 11940
rect 4169 11452 4477 11461
rect 4169 11450 4175 11452
rect 4231 11450 4255 11452
rect 4311 11450 4335 11452
rect 4391 11450 4415 11452
rect 4471 11450 4477 11452
rect 4231 11398 4233 11450
rect 4413 11398 4415 11450
rect 4169 11396 4175 11398
rect 4231 11396 4255 11398
rect 4311 11396 4335 11398
rect 4391 11396 4415 11398
rect 4471 11396 4477 11398
rect 4169 11387 4477 11396
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2884 9178 2912 9930
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2976 8974 3004 11018
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10742 3464 10950
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 7886 2176 8774
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 3528 7478 3556 11222
rect 5184 11218 5212 12310
rect 7392 12306 7420 13126
rect 7576 12986 7604 13466
rect 7668 13433 7696 14282
rect 7654 13424 7710 13433
rect 7654 13359 7710 13368
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7668 12238 7696 13359
rect 7760 13326 7788 14350
rect 7944 14006 7972 14350
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8220 14006 8248 14214
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7852 12850 7880 13670
rect 7944 13546 7972 13942
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 7944 13518 8064 13546
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12986 7972 13262
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8036 12850 8064 13518
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8128 12782 8156 13330
rect 8404 13326 8432 13874
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8312 12594 8340 13194
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8220 12566 8340 12594
rect 8220 12434 8248 12566
rect 8220 12406 8340 12434
rect 8312 12238 8340 12406
rect 8404 12374 8432 12786
rect 8496 12442 8524 14010
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8588 13462 8616 13874
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8680 12850 8708 14214
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8772 12782 8800 14282
rect 8864 13870 8892 14350
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13734 8892 13806
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8864 13462 8892 13670
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 8852 13320 8904 13326
rect 8850 13288 8852 13297
rect 8904 13288 8906 13297
rect 8850 13223 8906 13232
rect 9034 13288 9090 13297
rect 9034 13223 9090 13232
rect 8760 12776 8812 12782
rect 8864 12753 8892 13223
rect 8760 12718 8812 12724
rect 8850 12744 8906 12753
rect 9048 12714 9076 13223
rect 8850 12679 8906 12688
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9140 12646 9168 13738
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 9232 11354 9260 16730
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9324 13297 9352 14554
rect 9416 14414 9444 16662
rect 9692 15570 9720 19246
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9784 16658 9812 17206
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9876 16794 9904 17138
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9876 16250 9904 16526
rect 9968 16250 9996 20402
rect 10244 20330 10272 20878
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10336 20262 10364 20878
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10322 20088 10378 20097
rect 10322 20023 10378 20032
rect 10336 19394 10364 20023
rect 10428 19854 10456 22374
rect 10520 21962 10548 23122
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10704 22438 10732 23054
rect 10980 22642 11008 23462
rect 11072 23118 11100 24278
rect 11268 23964 11576 23973
rect 11268 23962 11274 23964
rect 11330 23962 11354 23964
rect 11410 23962 11434 23964
rect 11490 23962 11514 23964
rect 11570 23962 11576 23964
rect 11330 23910 11332 23962
rect 11512 23910 11514 23962
rect 11268 23908 11274 23910
rect 11330 23908 11354 23910
rect 11410 23908 11434 23910
rect 11490 23908 11514 23910
rect 11570 23908 11576 23910
rect 11268 23899 11576 23908
rect 11716 23730 11744 24822
rect 12268 24818 12296 25978
rect 12452 25906 12480 26182
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12360 25430 12388 25842
rect 12348 25424 12400 25430
rect 12348 25366 12400 25372
rect 12452 25294 12480 25842
rect 12728 25294 12756 26726
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12912 25770 12940 26318
rect 12900 25764 12952 25770
rect 12900 25706 12952 25712
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12452 25158 12480 25230
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12268 24682 12296 24754
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12452 24614 12480 25094
rect 12544 24750 12572 25230
rect 12808 24948 12860 24954
rect 12808 24890 12860 24896
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11152 23112 11204 23118
rect 11428 23112 11480 23118
rect 11152 23054 11204 23060
rect 11426 23080 11428 23089
rect 11704 23112 11756 23118
rect 11480 23080 11482 23089
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10608 22332 10916 22341
rect 10608 22330 10614 22332
rect 10670 22330 10694 22332
rect 10750 22330 10774 22332
rect 10830 22330 10854 22332
rect 10910 22330 10916 22332
rect 10670 22278 10672 22330
rect 10852 22278 10854 22330
rect 10608 22276 10614 22278
rect 10670 22276 10694 22278
rect 10750 22276 10774 22278
rect 10830 22276 10854 22278
rect 10910 22276 10916 22278
rect 10608 22267 10916 22276
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10612 21434 10640 22170
rect 11072 22137 11100 22510
rect 11164 22234 11192 23054
rect 11704 23054 11756 23060
rect 11426 23015 11482 23024
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11268 22876 11576 22885
rect 11268 22874 11274 22876
rect 11330 22874 11354 22876
rect 11410 22874 11434 22876
rect 11490 22874 11514 22876
rect 11570 22874 11576 22876
rect 11330 22822 11332 22874
rect 11512 22822 11514 22874
rect 11268 22820 11274 22822
rect 11330 22820 11354 22822
rect 11410 22820 11434 22822
rect 11490 22820 11514 22822
rect 11570 22820 11576 22822
rect 11268 22811 11576 22820
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11348 22234 11376 22374
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11058 22128 11114 22137
rect 11532 22098 11560 22714
rect 11624 22166 11652 22918
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11058 22063 11114 22072
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11612 22024 11664 22030
rect 11610 21992 11612 22001
rect 11664 21992 11666 22001
rect 11610 21927 11666 21936
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10520 21406 10640 21434
rect 10520 20398 10548 21406
rect 10608 21244 10916 21253
rect 10608 21242 10614 21244
rect 10670 21242 10694 21244
rect 10750 21242 10774 21244
rect 10830 21242 10854 21244
rect 10910 21242 10916 21244
rect 10670 21190 10672 21242
rect 10852 21190 10854 21242
rect 10608 21188 10614 21190
rect 10670 21188 10694 21190
rect 10750 21188 10774 21190
rect 10830 21188 10854 21190
rect 10910 21188 10916 21190
rect 10608 21179 10916 21188
rect 10980 20466 11008 21830
rect 11268 21788 11576 21797
rect 11268 21786 11274 21788
rect 11330 21786 11354 21788
rect 11410 21786 11434 21788
rect 11490 21786 11514 21788
rect 11570 21786 11576 21788
rect 11330 21734 11332 21786
rect 11512 21734 11514 21786
rect 11268 21732 11274 21734
rect 11330 21732 11354 21734
rect 11410 21732 11434 21734
rect 11490 21732 11514 21734
rect 11570 21732 11576 21734
rect 11268 21723 11576 21732
rect 11268 20700 11576 20709
rect 11268 20698 11274 20700
rect 11330 20698 11354 20700
rect 11410 20698 11434 20700
rect 11490 20698 11514 20700
rect 11570 20698 11576 20700
rect 11330 20646 11332 20698
rect 11512 20646 11514 20698
rect 11268 20644 11274 20646
rect 11330 20644 11354 20646
rect 11410 20644 11434 20646
rect 11490 20644 11514 20646
rect 11570 20644 11576 20646
rect 11268 20635 11576 20644
rect 11716 20602 11744 23054
rect 11808 22642 11836 23190
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11900 22778 11928 23054
rect 12084 22982 12112 23462
rect 12452 23322 12480 24550
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11992 22681 12020 22714
rect 11978 22672 12034 22681
rect 11796 22636 11848 22642
rect 11978 22607 12034 22616
rect 11796 22578 11848 22584
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10888 20346 10916 20402
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19514 10456 19790
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10414 19408 10470 19417
rect 10048 19372 10100 19378
rect 10336 19366 10414 19394
rect 10414 19343 10470 19352
rect 10048 19314 10100 19320
rect 10060 18766 10088 19314
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18970 10272 19178
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10048 18760 10100 18766
rect 10100 18720 10180 18748
rect 10048 18702 10100 18708
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 17882 10088 18566
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10152 17066 10180 18720
rect 10244 18426 10272 18906
rect 10428 18902 10456 19343
rect 10520 18970 10548 20334
rect 10888 20318 11008 20346
rect 10608 20156 10916 20165
rect 10608 20154 10614 20156
rect 10670 20154 10694 20156
rect 10750 20154 10774 20156
rect 10830 20154 10854 20156
rect 10910 20154 10916 20156
rect 10670 20102 10672 20154
rect 10852 20102 10854 20154
rect 10608 20100 10614 20102
rect 10670 20100 10694 20102
rect 10750 20100 10774 20102
rect 10830 20100 10854 20102
rect 10910 20100 10916 20102
rect 10608 20091 10916 20100
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10612 19378 10640 19450
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10888 19310 10916 19790
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10608 19068 10916 19077
rect 10608 19066 10614 19068
rect 10670 19066 10694 19068
rect 10750 19066 10774 19068
rect 10830 19066 10854 19068
rect 10910 19066 10916 19068
rect 10670 19014 10672 19066
rect 10852 19014 10854 19066
rect 10608 19012 10614 19014
rect 10670 19012 10694 19014
rect 10750 19012 10774 19014
rect 10830 19012 10854 19014
rect 10910 19012 10916 19014
rect 10608 19003 10916 19012
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10152 15910 10180 17002
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9310 13288 9366 13297
rect 9310 13223 9366 13232
rect 9416 12918 9444 14350
rect 9692 14074 9720 14350
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9784 13938 9812 14214
rect 10060 14006 10088 15506
rect 10244 14550 10272 18226
rect 10336 17678 10364 18226
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10520 17542 10548 18702
rect 10608 17980 10916 17989
rect 10608 17978 10614 17980
rect 10670 17978 10694 17980
rect 10750 17978 10774 17980
rect 10830 17978 10854 17980
rect 10910 17978 10916 17980
rect 10670 17926 10672 17978
rect 10852 17926 10854 17978
rect 10608 17924 10614 17926
rect 10670 17924 10694 17926
rect 10750 17924 10774 17926
rect 10830 17924 10854 17926
rect 10910 17924 10916 17926
rect 10608 17915 10916 17924
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10704 17610 10732 17750
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10612 17202 10640 17478
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10888 17134 10916 17750
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10520 15994 10548 17070
rect 10608 16892 10916 16901
rect 10608 16890 10614 16892
rect 10670 16890 10694 16892
rect 10750 16890 10774 16892
rect 10830 16890 10854 16892
rect 10910 16890 10916 16892
rect 10670 16838 10672 16890
rect 10852 16838 10854 16890
rect 10608 16836 10614 16838
rect 10670 16836 10694 16838
rect 10750 16836 10774 16838
rect 10830 16836 10854 16838
rect 10910 16836 10916 16838
rect 10608 16827 10916 16836
rect 10980 16454 11008 20318
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19922 11192 20198
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19378 11100 19654
rect 11164 19378 11192 19858
rect 11348 19854 11376 20470
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 20058 11836 20402
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19938 11836 19994
rect 11624 19922 11836 19938
rect 11612 19916 11836 19922
rect 11664 19910 11836 19916
rect 11612 19858 11664 19864
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11794 19816 11850 19825
rect 11612 19780 11664 19786
rect 11794 19751 11850 19760
rect 11612 19722 11664 19728
rect 11268 19612 11576 19621
rect 11268 19610 11274 19612
rect 11330 19610 11354 19612
rect 11410 19610 11434 19612
rect 11490 19610 11514 19612
rect 11570 19610 11576 19612
rect 11330 19558 11332 19610
rect 11512 19558 11514 19610
rect 11268 19556 11274 19558
rect 11330 19556 11354 19558
rect 11410 19556 11434 19558
rect 11490 19556 11514 19558
rect 11570 19556 11576 19558
rect 11268 19547 11576 19556
rect 11624 19514 11652 19722
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11808 19378 11836 19751
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18834 11100 19178
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11268 18524 11576 18533
rect 11268 18522 11274 18524
rect 11330 18522 11354 18524
rect 11410 18522 11434 18524
rect 11490 18522 11514 18524
rect 11570 18522 11576 18524
rect 11330 18470 11332 18522
rect 11512 18470 11514 18522
rect 11268 18468 11274 18470
rect 11330 18468 11354 18470
rect 11410 18468 11434 18470
rect 11490 18468 11514 18470
rect 11570 18468 11576 18470
rect 11268 18459 11576 18468
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11072 16998 11100 17818
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17338 11192 17478
rect 11268 17436 11576 17445
rect 11268 17434 11274 17436
rect 11330 17434 11354 17436
rect 11410 17434 11434 17436
rect 11490 17434 11514 17436
rect 11570 17434 11576 17436
rect 11330 17382 11332 17434
rect 11512 17382 11514 17434
rect 11268 17380 11274 17382
rect 11330 17380 11354 17382
rect 11410 17380 11434 17382
rect 11490 17380 11514 17382
rect 11570 17380 11576 17382
rect 11268 17371 11576 17380
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16522 11100 16934
rect 11164 16538 11192 17274
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11256 16794 11284 17002
rect 11624 16794 11652 17070
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11164 16522 11376 16538
rect 11060 16516 11112 16522
rect 11164 16516 11388 16522
rect 11164 16510 11336 16516
rect 11060 16458 11112 16464
rect 11336 16458 11388 16464
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 11268 16348 11576 16357
rect 11268 16346 11274 16348
rect 11330 16346 11354 16348
rect 11410 16346 11434 16348
rect 11490 16346 11514 16348
rect 11570 16346 11576 16348
rect 11330 16294 11332 16346
rect 11512 16294 11514 16346
rect 11268 16292 11274 16294
rect 11330 16292 11354 16294
rect 11410 16292 11434 16294
rect 11490 16292 11514 16294
rect 11570 16292 11576 16294
rect 11268 16283 11576 16292
rect 11334 16144 11390 16153
rect 11624 16114 11652 16594
rect 11716 16454 11744 19246
rect 11900 19242 11928 22374
rect 12084 22166 12112 22918
rect 12176 22556 12204 23122
rect 12636 23118 12664 23666
rect 12820 23322 12848 24890
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12912 24410 12940 24754
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 13004 24138 13032 25638
rect 13096 24818 13124 26726
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 13188 25498 13216 26250
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13372 25498 13400 25774
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13096 23798 13124 24550
rect 13188 24138 13216 24618
rect 13280 24410 13308 24754
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13084 23792 13136 23798
rect 13084 23734 13136 23740
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12440 22704 12492 22710
rect 12492 22664 12572 22692
rect 12440 22646 12492 22652
rect 12256 22568 12308 22574
rect 12176 22528 12256 22556
rect 12256 22510 12308 22516
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12268 22438 12296 22510
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12268 22030 12296 22374
rect 12452 22234 12480 22510
rect 12544 22234 12572 22664
rect 12728 22545 12756 22918
rect 12912 22642 12940 22918
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12714 22536 12770 22545
rect 13004 22506 13032 23190
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 12714 22471 12770 22480
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 13280 22438 13308 22986
rect 13372 22642 13400 25434
rect 13464 24818 13492 26386
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13556 25838 13584 26182
rect 13832 26042 13860 26182
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 14108 25702 14136 26318
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13556 24954 13584 25230
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13740 24206 13768 25298
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13556 23730 13584 24006
rect 13832 23866 13860 24822
rect 13924 24614 13952 25434
rect 14292 25294 14320 26318
rect 14384 25362 14412 26522
rect 14844 26382 14872 27066
rect 16212 26784 16264 26790
rect 16212 26726 16264 26732
rect 15844 26512 15896 26518
rect 15844 26454 15896 26460
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14476 25498 14504 26318
rect 14740 26240 14792 26246
rect 14740 26182 14792 26188
rect 14752 25974 14780 26182
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14476 25294 14504 25434
rect 14568 25294 14596 25638
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24750 14136 25094
rect 14476 24886 14504 25230
rect 14568 24954 14596 25230
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 14844 23730 14872 26318
rect 15764 26246 15792 26386
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 25906 15792 26182
rect 15856 25974 15884 26454
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15844 25968 15896 25974
rect 15844 25910 15896 25916
rect 16040 25906 16068 26318
rect 16224 26314 16252 26726
rect 16212 26308 16264 26314
rect 16212 26250 16264 26256
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 15120 24750 15148 25162
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 13832 23526 13860 23666
rect 15212 23662 15240 25230
rect 15660 25220 15712 25226
rect 15660 25162 15712 25168
rect 15672 24886 15700 25162
rect 15764 25158 15792 25842
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15948 24886 15976 25842
rect 16040 25498 16068 25842
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 16224 25294 16252 26250
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 16396 25220 16448 25226
rect 16396 25162 16448 25168
rect 16408 24954 16436 25162
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 13832 23118 13860 23462
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22778 13492 22918
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12452 21622 12480 22170
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 13280 21350 13308 22170
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13464 21010 13492 22714
rect 13832 22642 13860 23054
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 14200 22574 14228 23122
rect 14384 22710 14412 23462
rect 15212 22778 15240 23598
rect 15672 23322 15700 24822
rect 15948 24410 15976 24822
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15842 23216 15898 23225
rect 15842 23151 15898 23160
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 15856 22642 15884 23151
rect 16316 23050 16344 23462
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16592 22658 16620 27338
rect 17707 27228 18015 27237
rect 17707 27226 17713 27228
rect 17769 27226 17793 27228
rect 17849 27226 17873 27228
rect 17929 27226 17953 27228
rect 18009 27226 18015 27228
rect 17769 27174 17771 27226
rect 17951 27174 17953 27226
rect 17707 27172 17713 27174
rect 17769 27172 17793 27174
rect 17849 27172 17873 27174
rect 17929 27172 17953 27174
rect 18009 27172 18015 27174
rect 17707 27163 18015 27172
rect 24146 27228 24454 27237
rect 24146 27226 24152 27228
rect 24208 27226 24232 27228
rect 24288 27226 24312 27228
rect 24368 27226 24392 27228
rect 24448 27226 24454 27228
rect 24208 27174 24210 27226
rect 24390 27174 24392 27226
rect 24146 27172 24152 27174
rect 24208 27172 24232 27174
rect 24288 27172 24312 27174
rect 24368 27172 24392 27174
rect 24448 27172 24454 27174
rect 24146 27163 24454 27172
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16684 25838 16712 26386
rect 16868 26314 16896 26726
rect 17047 26684 17355 26693
rect 17047 26682 17053 26684
rect 17109 26682 17133 26684
rect 17189 26682 17213 26684
rect 17269 26682 17293 26684
rect 17349 26682 17355 26684
rect 17109 26630 17111 26682
rect 17291 26630 17293 26682
rect 17047 26628 17053 26630
rect 17109 26628 17133 26630
rect 17189 26628 17213 26630
rect 17269 26628 17293 26630
rect 17349 26628 17355 26630
rect 17047 26619 17355 26628
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16684 25430 16712 25774
rect 17420 25702 17448 26318
rect 17512 26042 17540 26862
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 17707 26140 18015 26149
rect 17707 26138 17713 26140
rect 17769 26138 17793 26140
rect 17849 26138 17873 26140
rect 17929 26138 17953 26140
rect 18009 26138 18015 26140
rect 17769 26086 17771 26138
rect 17951 26086 17953 26138
rect 17707 26084 17713 26086
rect 17769 26084 17793 26086
rect 17849 26084 17873 26086
rect 17929 26084 17953 26086
rect 18009 26084 18015 26086
rect 17707 26075 18015 26084
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 18064 25974 18092 26182
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17047 25596 17355 25605
rect 17047 25594 17053 25596
rect 17109 25594 17133 25596
rect 17189 25594 17213 25596
rect 17269 25594 17293 25596
rect 17349 25594 17355 25596
rect 17109 25542 17111 25594
rect 17291 25542 17293 25594
rect 17047 25540 17053 25542
rect 17109 25540 17133 25542
rect 17189 25540 17213 25542
rect 17269 25540 17293 25542
rect 17349 25540 17355 25542
rect 17047 25531 17355 25540
rect 16672 25424 16724 25430
rect 16672 25366 16724 25372
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 16500 22630 16620 22658
rect 16684 22642 16712 23122
rect 16868 23118 16896 25094
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16960 22778 16988 25366
rect 17707 25052 18015 25061
rect 17707 25050 17713 25052
rect 17769 25050 17793 25052
rect 17849 25050 17873 25052
rect 17929 25050 17953 25052
rect 18009 25050 18015 25052
rect 17769 24998 17771 25050
rect 17951 24998 17953 25050
rect 17707 24996 17713 24998
rect 17769 24996 17793 24998
rect 17849 24996 17873 24998
rect 17929 24996 17953 24998
rect 18009 24996 18015 24998
rect 17707 24987 18015 24996
rect 18156 24800 18184 26726
rect 18984 26586 19012 26998
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 18972 26580 19024 26586
rect 18972 26522 19024 26528
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 19352 25906 19380 26182
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18236 24812 18288 24818
rect 18156 24772 18236 24800
rect 18236 24754 18288 24760
rect 17047 24508 17355 24517
rect 17047 24506 17053 24508
rect 17109 24506 17133 24508
rect 17189 24506 17213 24508
rect 17269 24506 17293 24508
rect 17349 24506 17355 24508
rect 17109 24454 17111 24506
rect 17291 24454 17293 24506
rect 17047 24452 17053 24454
rect 17109 24452 17133 24454
rect 17189 24452 17213 24454
rect 17269 24452 17293 24454
rect 17349 24452 17355 24454
rect 17047 24443 17355 24452
rect 17707 23964 18015 23973
rect 17707 23962 17713 23964
rect 17769 23962 17793 23964
rect 17849 23962 17873 23964
rect 17929 23962 17953 23964
rect 18009 23962 18015 23964
rect 17769 23910 17771 23962
rect 17951 23910 17953 23962
rect 17707 23908 17713 23910
rect 17769 23908 17793 23910
rect 17849 23908 17873 23910
rect 17929 23908 17953 23910
rect 18009 23908 18015 23910
rect 17707 23899 18015 23908
rect 18248 23798 18276 24754
rect 18524 24614 18552 25366
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18616 24818 18644 25162
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18800 24818 18828 25094
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19064 24812 19116 24818
rect 19116 24772 19288 24800
rect 19064 24754 19116 24760
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 24274 18552 24550
rect 18616 24342 18644 24754
rect 18984 24410 19012 24754
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19260 24562 19288 24772
rect 19352 24682 19380 25230
rect 19444 24818 19472 26250
rect 19628 26042 19656 26250
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 19720 25498 19748 26862
rect 19996 26450 20024 26862
rect 23486 26684 23794 26693
rect 23486 26682 23492 26684
rect 23548 26682 23572 26684
rect 23628 26682 23652 26684
rect 23708 26682 23732 26684
rect 23788 26682 23794 26684
rect 23548 26630 23550 26682
rect 23730 26630 23732 26682
rect 23486 26628 23492 26630
rect 23548 26628 23572 26630
rect 23628 26628 23652 26630
rect 23708 26628 23732 26630
rect 23788 26628 23794 26630
rect 23486 26619 23794 26628
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 19536 24562 19564 25230
rect 19628 24886 19656 25230
rect 19616 24880 19668 24886
rect 19616 24822 19668 24828
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 17047 23420 17355 23429
rect 17047 23418 17053 23420
rect 17109 23418 17133 23420
rect 17189 23418 17213 23420
rect 17269 23418 17293 23420
rect 17349 23418 17355 23420
rect 17109 23366 17111 23418
rect 17291 23366 17293 23418
rect 17047 23364 17053 23366
rect 17109 23364 17133 23366
rect 17189 23364 17213 23366
rect 17269 23364 17293 23366
rect 17349 23364 17355 23366
rect 17047 23355 17355 23364
rect 18248 23089 18276 23734
rect 18524 23118 18552 24210
rect 19168 24206 19196 24550
rect 19260 24534 19564 24562
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23798 19196 24142
rect 19260 24138 19288 24534
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19260 23118 19288 24074
rect 19352 23730 19380 24278
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 19352 23254 19380 23530
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 18328 23112 18380 23118
rect 18234 23080 18290 23089
rect 18328 23054 18380 23060
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19248 23112 19300 23118
rect 19444 23100 19472 24346
rect 19812 23866 19840 24686
rect 19800 23860 19852 23866
rect 19628 23820 19800 23848
rect 19524 23112 19576 23118
rect 19444 23072 19524 23100
rect 19248 23054 19300 23060
rect 19524 23054 19576 23060
rect 18234 23015 18290 23024
rect 17707 22876 18015 22885
rect 17707 22874 17713 22876
rect 17769 22874 17793 22876
rect 17849 22874 17873 22876
rect 17929 22874 17953 22876
rect 18009 22874 18015 22876
rect 17769 22822 17771 22874
rect 17951 22822 17953 22874
rect 17707 22820 17713 22822
rect 17769 22820 17793 22822
rect 17849 22820 17873 22822
rect 17929 22820 17953 22822
rect 18009 22820 18015 22822
rect 17707 22811 18015 22820
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16672 22636 16724 22642
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14200 22234 14228 22510
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14660 21690 14688 22374
rect 16500 22114 16528 22630
rect 16672 22578 16724 22584
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16592 22234 16620 22510
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16396 22092 16448 22098
rect 16500 22086 16620 22114
rect 16396 22034 16448 22040
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15660 21956 15712 21962
rect 15660 21898 15712 21904
rect 15212 21690 15240 21898
rect 15672 21690 15700 21898
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15948 21622 15976 21966
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 13556 21078 13584 21558
rect 16408 21554 16436 22034
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 14016 21146 14044 21422
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 14476 20874 14504 21490
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14568 20777 14596 21422
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14554 20768 14610 20777
rect 14554 20703 14610 20712
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 12254 19952 12310 19961
rect 14476 19922 14504 20266
rect 12254 19887 12310 19896
rect 14464 19916 14516 19922
rect 12268 19854 12296 19887
rect 14464 19858 14516 19864
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 12544 18970 12572 19314
rect 12820 19174 12848 19722
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19446 13768 19654
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12820 18766 12848 19110
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12544 17678 12572 18158
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17882 12756 18090
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11334 16079 11336 16088
rect 11388 16079 11390 16088
rect 11612 16108 11664 16114
rect 11336 16050 11388 16056
rect 11612 16050 11664 16056
rect 10520 15966 11008 15994
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15434 10548 15846
rect 10608 15804 10916 15813
rect 10608 15802 10614 15804
rect 10670 15802 10694 15804
rect 10750 15802 10774 15804
rect 10830 15802 10854 15804
rect 10910 15802 10916 15804
rect 10670 15750 10672 15802
rect 10852 15750 10854 15802
rect 10608 15748 10614 15750
rect 10670 15748 10694 15750
rect 10750 15748 10774 15750
rect 10830 15748 10854 15750
rect 10910 15748 10916 15750
rect 10608 15739 10916 15748
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10608 14716 10916 14725
rect 10608 14714 10614 14716
rect 10670 14714 10694 14716
rect 10750 14714 10774 14716
rect 10830 14714 10854 14716
rect 10910 14714 10916 14716
rect 10670 14662 10672 14714
rect 10852 14662 10854 14714
rect 10608 14660 10614 14662
rect 10670 14660 10694 14662
rect 10750 14660 10774 14662
rect 10830 14660 10854 14662
rect 10910 14660 10916 14662
rect 10608 14651 10916 14660
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13326 10088 13670
rect 10608 13628 10916 13637
rect 10608 13626 10614 13628
rect 10670 13626 10694 13628
rect 10750 13626 10774 13628
rect 10830 13626 10854 13628
rect 10910 13626 10916 13628
rect 10670 13574 10672 13626
rect 10852 13574 10854 13626
rect 10608 13572 10614 13574
rect 10670 13572 10694 13574
rect 10750 13572 10774 13574
rect 10830 13572 10854 13574
rect 10910 13572 10916 13574
rect 10608 13563 10916 13572
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9600 12170 9628 12718
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 4080 11121 4108 11154
rect 4066 11112 4122 11121
rect 3884 11076 3936 11082
rect 4066 11047 4122 11056
rect 5356 11076 5408 11082
rect 3884 11018 3936 11024
rect 5356 11018 5408 11024
rect 3896 10674 3924 11018
rect 4829 10908 5137 10917
rect 4829 10906 4835 10908
rect 4891 10906 4915 10908
rect 4971 10906 4995 10908
rect 5051 10906 5075 10908
rect 5131 10906 5137 10908
rect 4891 10854 4893 10906
rect 5073 10854 5075 10906
rect 4829 10852 4835 10854
rect 4891 10852 4915 10854
rect 4971 10852 4995 10854
rect 5051 10852 5075 10854
rect 5131 10852 5137 10854
rect 4829 10843 5137 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4264 10674 4292 10746
rect 5276 10674 5304 10746
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 9654 3740 10406
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3988 9382 4016 10610
rect 4620 10600 4672 10606
rect 4540 10548 4620 10554
rect 4540 10542 4672 10548
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4540 10526 4660 10542
rect 4712 10532 4764 10538
rect 4080 10266 4108 10474
rect 4169 10364 4477 10373
rect 4169 10362 4175 10364
rect 4231 10362 4255 10364
rect 4311 10362 4335 10364
rect 4391 10362 4415 10364
rect 4471 10362 4477 10364
rect 4231 10310 4233 10362
rect 4413 10310 4415 10362
rect 4169 10308 4175 10310
rect 4231 10308 4255 10310
rect 4311 10308 4335 10310
rect 4391 10308 4415 10310
rect 4471 10308 4477 10310
rect 4169 10299 4477 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 9674 4108 10202
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4264 9722 4292 9930
rect 4252 9716 4304 9722
rect 4080 9646 4200 9674
rect 4252 9658 4304 9664
rect 3976 9376 4028 9382
rect 4172 9364 4200 9646
rect 4356 9518 4384 9930
rect 4540 9654 4568 10526
rect 4712 10474 4764 10480
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10198 4660 10406
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 3976 9318 4028 9324
rect 4080 9336 4200 9364
rect 4080 9042 4108 9336
rect 4169 9276 4477 9285
rect 4169 9274 4175 9276
rect 4231 9274 4255 9276
rect 4311 9274 4335 9276
rect 4391 9274 4415 9276
rect 4471 9274 4477 9276
rect 4231 9222 4233 9274
rect 4413 9222 4415 9274
rect 4169 9220 4175 9222
rect 4231 9220 4255 9222
rect 4311 9220 4335 9222
rect 4391 9220 4415 9222
rect 4471 9220 4477 9222
rect 4169 9211 4477 9220
rect 4632 9110 4660 9998
rect 4724 9586 4752 10474
rect 4804 10056 4856 10062
rect 4802 10024 4804 10033
rect 4908 10044 4936 10610
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10266 5120 10474
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5092 10130 5120 10202
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5184 10062 5212 10406
rect 5276 10130 5304 10610
rect 5368 10538 5396 11018
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 4988 10056 5040 10062
rect 4856 10024 4858 10033
rect 4908 10016 4988 10044
rect 4988 9998 5040 10004
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 4802 9959 4858 9968
rect 5000 9926 5028 9998
rect 4988 9920 5040 9926
rect 5040 9880 5212 9908
rect 4988 9862 5040 9868
rect 4829 9820 5137 9829
rect 4829 9818 4835 9820
rect 4891 9818 4915 9820
rect 4971 9818 4995 9820
rect 5051 9818 5075 9820
rect 5131 9818 5137 9820
rect 4891 9766 4893 9818
rect 5073 9766 5075 9818
rect 4829 9764 4835 9766
rect 4891 9764 4915 9766
rect 4971 9764 4995 9766
rect 5051 9764 5075 9766
rect 5131 9764 5137 9766
rect 4829 9755 5137 9764
rect 5184 9586 5212 9880
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5276 9382 5304 10066
rect 5354 10024 5410 10033
rect 5354 9959 5410 9968
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5368 9364 5396 9959
rect 5460 9636 5488 11154
rect 6734 11112 6790 11121
rect 6460 11076 6512 11082
rect 6734 11047 6790 11056
rect 6460 11018 6512 11024
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5552 10266 5580 10678
rect 6380 10674 6408 10950
rect 6472 10810 6500 11018
rect 6748 11014 6776 11047
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5644 10266 5672 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5816 10192 5868 10198
rect 5552 10140 5816 10146
rect 5552 10134 5868 10140
rect 5552 10118 5856 10134
rect 5552 10062 5580 10118
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5828 9722 5856 10118
rect 5920 10062 5948 10610
rect 6840 10198 6868 10678
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6840 10062 6868 10134
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5460 9608 5580 9636
rect 5448 9376 5500 9382
rect 5368 9336 5448 9364
rect 5184 9194 5212 9318
rect 5368 9194 5396 9336
rect 5448 9318 5500 9324
rect 5184 9166 5396 9194
rect 5460 9110 5488 9318
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4829 8732 5137 8741
rect 4829 8730 4835 8732
rect 4891 8730 4915 8732
rect 4971 8730 4995 8732
rect 5051 8730 5075 8732
rect 5131 8730 5137 8732
rect 4891 8678 4893 8730
rect 5073 8678 5075 8730
rect 4829 8676 4835 8678
rect 4891 8676 4915 8678
rect 4971 8676 4995 8678
rect 5051 8676 5075 8678
rect 5131 8676 5137 8678
rect 4829 8667 5137 8676
rect 5552 8498 5580 9608
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9364 5856 9522
rect 6012 9518 6040 9862
rect 6380 9722 6408 9930
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5908 9376 5960 9382
rect 5828 9336 5908 9364
rect 5908 9318 5960 9324
rect 5920 9042 5948 9318
rect 6012 9178 6040 9454
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6104 8974 6132 9318
rect 6196 9110 6224 9590
rect 6472 9586 6500 9930
rect 6932 9654 6960 10542
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9382 7052 9522
rect 7392 9518 7420 10610
rect 7484 10062 7512 10610
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 10062 7788 10202
rect 7852 10062 7880 10406
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7484 9586 7512 9998
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7576 9518 7604 9930
rect 7760 9586 7788 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7852 9654 7880 9862
rect 7944 9654 7972 9862
rect 8036 9722 8064 10746
rect 8128 10674 8156 10746
rect 8588 10674 8616 11154
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 8772 10810 8800 10950
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8680 10674 8708 10746
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8588 10538 8616 10610
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8220 10062 8248 10474
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10198 8524 10406
rect 8588 10198 8616 10474
rect 8680 10470 8708 10610
rect 9416 10606 9444 10678
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 8404 9586 8432 9862
rect 8588 9586 8616 10134
rect 8680 9586 8708 10406
rect 8772 10266 8800 10474
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8956 10062 8984 10542
rect 9048 10130 9076 10542
rect 9416 10146 9444 10542
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9324 10118 9444 10146
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9926 8984 9998
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9586 8984 9862
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7116 9178 7144 9454
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6196 8634 6224 9046
rect 8588 8838 8616 9522
rect 8680 9042 8708 9522
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 4169 8188 4477 8197
rect 4169 8186 4175 8188
rect 4231 8186 4255 8188
rect 4311 8186 4335 8188
rect 4391 8186 4415 8188
rect 4471 8186 4477 8188
rect 4231 8134 4233 8186
rect 4413 8134 4415 8186
rect 4169 8132 4175 8134
rect 4231 8132 4255 8134
rect 4311 8132 4335 8134
rect 4391 8132 4415 8134
rect 4471 8132 4477 8134
rect 4169 8123 4477 8132
rect 5552 8090 5580 8434
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3516 7472 3568 7478
rect 3516 7414 3568 7420
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6730 3096 7142
rect 3252 6866 3280 7210
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5642 2268 6054
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 2650 2452 5170
rect 3712 4146 3740 6734
rect 3804 6254 3832 7686
rect 3884 7336 3936 7342
rect 4172 7290 4200 7822
rect 4264 7546 4292 7822
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3884 7278 3936 7284
rect 3896 6798 3924 7278
rect 4080 7262 4200 7290
rect 4080 6882 4108 7262
rect 4169 7100 4477 7109
rect 4169 7098 4175 7100
rect 4231 7098 4255 7100
rect 4311 7098 4335 7100
rect 4391 7098 4415 7100
rect 4471 7098 4477 7100
rect 4231 7046 4233 7098
rect 4413 7046 4415 7098
rect 4169 7044 4175 7046
rect 4231 7044 4255 7046
rect 4311 7044 4335 7046
rect 4391 7044 4415 7046
rect 4471 7044 4477 7046
rect 4169 7035 4477 7044
rect 4080 6854 4476 6882
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4448 6730 4476 6854
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6390 3924 6598
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 4172 6322 4200 6666
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3792 6248 3844 6254
rect 4172 6202 4200 6258
rect 4448 6254 4476 6666
rect 4540 6458 4568 7822
rect 4829 7644 5137 7653
rect 4829 7642 4835 7644
rect 4891 7642 4915 7644
rect 4971 7642 4995 7644
rect 5051 7642 5075 7644
rect 5131 7642 5137 7644
rect 4891 7590 4893 7642
rect 5073 7590 5075 7642
rect 4829 7588 4835 7590
rect 4891 7588 4915 7590
rect 4971 7588 4995 7590
rect 5051 7588 5075 7590
rect 5131 7588 5137 7590
rect 4829 7579 5137 7588
rect 5644 7478 5672 7890
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4632 6322 4660 7346
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4816 6798 4844 7142
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 3792 6190 3844 6196
rect 4080 6174 4200 6202
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3712 3534 3740 4082
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3988 2990 4016 3878
rect 4080 3602 4108 6174
rect 4169 6012 4477 6021
rect 4169 6010 4175 6012
rect 4231 6010 4255 6012
rect 4311 6010 4335 6012
rect 4391 6010 4415 6012
rect 4471 6010 4477 6012
rect 4231 5958 4233 6010
rect 4413 5958 4415 6010
rect 4169 5956 4175 5958
rect 4231 5956 4255 5958
rect 4311 5956 4335 5958
rect 4391 5956 4415 5958
rect 4471 5956 4477 5958
rect 4169 5947 4477 5956
rect 4632 5914 4660 6258
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4169 4924 4477 4933
rect 4169 4922 4175 4924
rect 4231 4922 4255 4924
rect 4311 4922 4335 4924
rect 4391 4922 4415 4924
rect 4471 4922 4477 4924
rect 4231 4870 4233 4922
rect 4413 4870 4415 4922
rect 4169 4868 4175 4870
rect 4231 4868 4255 4870
rect 4311 4868 4335 4870
rect 4391 4868 4415 4870
rect 4471 4868 4477 4870
rect 4169 4859 4477 4868
rect 4724 4622 4752 6666
rect 4829 6556 5137 6565
rect 4829 6554 4835 6556
rect 4891 6554 4915 6556
rect 4971 6554 4995 6556
rect 5051 6554 5075 6556
rect 5131 6554 5137 6556
rect 4891 6502 4893 6554
rect 5073 6502 5075 6554
rect 4829 6500 4835 6502
rect 4891 6500 4915 6502
rect 4971 6500 4995 6502
rect 5051 6500 5075 6502
rect 5131 6500 5137 6502
rect 4829 6491 5137 6500
rect 5184 6458 5212 7278
rect 5368 7018 5396 7346
rect 5368 7002 5488 7018
rect 5368 6996 5500 7002
rect 5368 6990 5448 6996
rect 5368 6798 5396 6990
rect 5448 6938 5500 6944
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4816 6322 4844 6394
rect 5276 6322 5304 6734
rect 5460 6390 5488 6802
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5276 5914 5304 6258
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5778 5396 6258
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 4829 5468 5137 5477
rect 4829 5466 4835 5468
rect 4891 5466 4915 5468
rect 4971 5466 4995 5468
rect 5051 5466 5075 5468
rect 5131 5466 5137 5468
rect 4891 5414 4893 5466
rect 5073 5414 5075 5466
rect 4829 5412 4835 5414
rect 4891 5412 4915 5414
rect 4971 5412 4995 5414
rect 5051 5412 5075 5414
rect 5131 5412 5137 5414
rect 4829 5403 5137 5412
rect 5184 4622 5212 5714
rect 5460 5642 5488 6326
rect 5644 5710 5672 7414
rect 7208 7410 7236 7822
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7484 7546 7512 7754
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 5736 6322 5764 7346
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 6798 5948 7142
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5920 6390 5948 6598
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6012 6322 6040 6598
rect 6104 6458 6132 6734
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5736 6186 5764 6258
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5644 5370 5672 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4282 4292 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4172 3942 4200 4150
rect 4448 4146 4476 4490
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4169 3836 4477 3845
rect 4169 3834 4175 3836
rect 4231 3834 4255 3836
rect 4311 3834 4335 3836
rect 4391 3834 4415 3836
rect 4471 3834 4477 3836
rect 4231 3782 4233 3834
rect 4413 3782 4415 3834
rect 4169 3780 4175 3782
rect 4231 3780 4255 3782
rect 4311 3780 4335 3782
rect 4391 3780 4415 3782
rect 4471 3780 4477 3782
rect 4169 3771 4477 3780
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3126 4108 3538
rect 4252 3528 4304 3534
rect 4540 3516 4568 4422
rect 4724 4078 4752 4558
rect 4829 4380 5137 4389
rect 4829 4378 4835 4380
rect 4891 4378 4915 4380
rect 4971 4378 4995 4380
rect 5051 4378 5075 4380
rect 5131 4378 5137 4380
rect 4891 4326 4893 4378
rect 5073 4326 5075 4378
rect 4829 4324 4835 4326
rect 4891 4324 4915 4326
rect 4971 4324 4995 4326
rect 5051 4324 5075 4326
rect 5131 4324 5137 4326
rect 4829 4315 5137 4324
rect 5184 4214 5212 4558
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4304 3488 4568 3516
rect 4252 3470 4304 3476
rect 4632 3126 4660 3946
rect 4829 3292 5137 3301
rect 4829 3290 4835 3292
rect 4891 3290 4915 3292
rect 4971 3290 4995 3292
rect 5051 3290 5075 3292
rect 5131 3290 5137 3292
rect 4891 3238 4893 3290
rect 5073 3238 5075 3290
rect 4829 3236 4835 3238
rect 4891 3236 4915 3238
rect 4971 3236 4995 3238
rect 5051 3236 5075 3238
rect 5131 3236 5137 3238
rect 4829 3227 5137 3236
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 5552 2922 5580 4490
rect 5736 4146 5764 6122
rect 6012 5642 6040 6122
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6012 5030 6040 5578
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5736 3738 5764 4082
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5736 3534 5764 3674
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5828 2990 5856 4082
rect 6012 3194 6040 4966
rect 6196 4690 6224 6054
rect 6288 5914 6316 6734
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 6118 6684 6190
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5930 6684 6054
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6564 5902 6684 5930
rect 6564 5846 6592 5902
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6288 4554 6316 5306
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 3942 6316 4490
rect 6380 4214 6408 4558
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6196 3126 6224 3878
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6288 2990 6316 3878
rect 6380 3602 6408 4150
rect 6564 4146 6592 5782
rect 6748 5710 6776 6258
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5778 6960 6190
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 4146 6776 5646
rect 6932 5302 6960 5714
rect 7208 5574 7236 7346
rect 8220 7342 8248 7754
rect 8312 7410 8340 7822
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 6322 7328 7210
rect 8220 7002 8248 7278
rect 8312 7002 8340 7346
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8220 6390 8248 6938
rect 8404 6798 8432 8298
rect 8680 7274 8708 8978
rect 9048 8498 9076 10066
rect 9324 10062 9352 10118
rect 9508 10062 9536 10202
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9324 9654 9352 9998
rect 9968 9994 9996 10950
rect 10336 10130 10364 13262
rect 10608 12540 10916 12549
rect 10608 12538 10614 12540
rect 10670 12538 10694 12540
rect 10750 12538 10774 12540
rect 10830 12538 10854 12540
rect 10910 12538 10916 12540
rect 10670 12486 10672 12538
rect 10852 12486 10854 12538
rect 10608 12484 10614 12486
rect 10670 12484 10694 12486
rect 10750 12484 10774 12486
rect 10830 12484 10854 12486
rect 10910 12484 10916 12486
rect 10608 12475 10916 12484
rect 10980 12434 11008 15966
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15434 11284 15846
rect 11624 15706 11652 16050
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11268 15260 11576 15269
rect 11268 15258 11274 15260
rect 11330 15258 11354 15260
rect 11410 15258 11434 15260
rect 11490 15258 11514 15260
rect 11570 15258 11576 15260
rect 11330 15206 11332 15258
rect 11512 15206 11514 15258
rect 11268 15204 11274 15206
rect 11330 15204 11354 15206
rect 11410 15204 11434 15206
rect 11490 15204 11514 15206
rect 11570 15204 11576 15206
rect 11268 15195 11576 15204
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11268 14172 11576 14181
rect 11268 14170 11274 14172
rect 11330 14170 11354 14172
rect 11410 14170 11434 14172
rect 11490 14170 11514 14172
rect 11570 14170 11576 14172
rect 11330 14118 11332 14170
rect 11512 14118 11514 14170
rect 11268 14116 11274 14118
rect 11330 14116 11354 14118
rect 11410 14116 11434 14118
rect 11490 14116 11514 14118
rect 11570 14116 11576 14118
rect 11268 14107 11576 14116
rect 11716 13938 11744 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11072 12918 11100 13670
rect 11164 13258 11192 13670
rect 11624 13512 11652 13874
rect 11624 13484 11744 13512
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11268 13084 11576 13093
rect 11268 13082 11274 13084
rect 11330 13082 11354 13084
rect 11410 13082 11434 13084
rect 11490 13082 11514 13084
rect 11570 13082 11576 13084
rect 11330 13030 11332 13082
rect 11512 13030 11514 13082
rect 11268 13028 11274 13030
rect 11330 13028 11354 13030
rect 11410 13028 11434 13030
rect 11490 13028 11514 13030
rect 11570 13028 11576 13030
rect 11268 13019 11576 13028
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11440 12442 11468 12922
rect 11624 12850 11652 13330
rect 11716 12986 11744 13484
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 10520 12406 11008 12434
rect 11428 12436 11480 12442
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 10428 9654 10456 10610
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9140 7886 9168 8502
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7478 8800 7686
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8772 7002 8800 7414
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8956 6798 8984 7346
rect 9140 7313 9168 7346
rect 9220 7336 9272 7342
rect 9126 7304 9182 7313
rect 9220 7278 9272 7284
rect 9126 7239 9182 7248
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 6866 9168 7142
rect 9232 7002 9260 7278
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9600 6905 9628 7890
rect 9784 7818 9812 8230
rect 10152 7886 10180 8842
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 10152 7342 10180 7822
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10322 7304 10378 7313
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9586 6896 9642 6905
rect 9128 6860 9180 6866
rect 9586 6831 9642 6840
rect 9680 6860 9732 6866
rect 9128 6802 9180 6808
rect 8392 6792 8444 6798
rect 8484 6792 8536 6798
rect 8392 6734 8444 6740
rect 8482 6760 8484 6769
rect 8944 6792 8996 6798
rect 8536 6760 8538 6769
rect 8944 6734 8996 6740
rect 8482 6695 8538 6704
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8496 6322 8524 6598
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9128 6384 9180 6390
rect 8942 6352 8998 6361
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 8484 6316 8536 6322
rect 9128 6326 9180 6332
rect 8942 6287 8944 6296
rect 8484 6258 8536 6264
rect 8996 6287 8998 6296
rect 8944 6258 8996 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 6118 7512 6190
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 8128 4826 8156 6054
rect 8956 5710 8984 6258
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 9140 5234 9168 6326
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5642 9260 6190
rect 9508 5710 9536 6394
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9232 5166 9260 5578
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9508 5234 9536 5510
rect 9600 5302 9628 6831
rect 9680 6802 9732 6808
rect 9692 6633 9720 6802
rect 9784 6798 9812 7142
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9678 6624 9734 6633
rect 9678 6559 9734 6568
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9680 6384 9732 6390
rect 9968 6361 9996 6394
rect 9680 6326 9732 6332
rect 9954 6352 10010 6361
rect 9692 5914 9720 6326
rect 9954 6287 10010 6296
rect 9772 6248 9824 6254
rect 9824 6208 9904 6236
rect 9772 6190 9824 6196
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9784 5642 9812 6054
rect 9876 5846 9904 6208
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8312 4690 8340 4966
rect 10060 4826 10088 7278
rect 10322 7239 10378 7248
rect 10336 7002 10364 7239
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6633 10272 6734
rect 10230 6624 10286 6633
rect 10230 6559 10286 6568
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10152 5914 10180 6190
rect 10244 6118 10272 6559
rect 10428 6254 10456 6938
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10520 5794 10548 12406
rect 11808 12434 11836 16934
rect 12360 16590 12388 17614
rect 12820 16998 12848 18702
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13556 18086 13584 18158
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17882 13584 18022
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13740 17678 13768 18226
rect 14200 18222 14228 19110
rect 14568 18426 14596 19314
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13174 17232 13230 17241
rect 13174 17167 13230 17176
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 11900 16250 11928 16390
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15570 12112 15982
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 14006 12112 15506
rect 12268 14346 12296 16390
rect 12360 16182 12388 16390
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 15706 12388 15982
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12084 13394 12112 13942
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12176 12986 12204 13806
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11428 12378 11480 12384
rect 11624 12406 11836 12434
rect 11268 11996 11576 12005
rect 11268 11994 11274 11996
rect 11330 11994 11354 11996
rect 11410 11994 11434 11996
rect 11490 11994 11514 11996
rect 11570 11994 11576 11996
rect 11330 11942 11332 11994
rect 11512 11942 11514 11994
rect 11268 11940 11274 11942
rect 11330 11940 11354 11942
rect 11410 11940 11434 11942
rect 11490 11940 11514 11942
rect 11570 11940 11576 11942
rect 11268 11931 11576 11940
rect 10608 11452 10916 11461
rect 10608 11450 10614 11452
rect 10670 11450 10694 11452
rect 10750 11450 10774 11452
rect 10830 11450 10854 11452
rect 10910 11450 10916 11452
rect 10670 11398 10672 11450
rect 10852 11398 10854 11450
rect 10608 11396 10614 11398
rect 10670 11396 10694 11398
rect 10750 11396 10774 11398
rect 10830 11396 10854 11398
rect 10910 11396 10916 11398
rect 10608 11387 10916 11396
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10656 11100 11018
rect 11164 10810 11192 11086
rect 11268 10908 11576 10917
rect 11268 10906 11274 10908
rect 11330 10906 11354 10908
rect 11410 10906 11434 10908
rect 11490 10906 11514 10908
rect 11570 10906 11576 10908
rect 11330 10854 11332 10906
rect 11512 10854 11514 10906
rect 11268 10852 11274 10854
rect 11330 10852 11354 10854
rect 11410 10852 11434 10854
rect 11490 10852 11514 10854
rect 11570 10852 11576 10854
rect 11268 10843 11576 10852
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11152 10668 11204 10674
rect 11072 10628 11152 10656
rect 11152 10610 11204 10616
rect 10608 10364 10916 10373
rect 10608 10362 10614 10364
rect 10670 10362 10694 10364
rect 10750 10362 10774 10364
rect 10830 10362 10854 10364
rect 10910 10362 10916 10364
rect 10670 10310 10672 10362
rect 10852 10310 10854 10362
rect 10608 10308 10614 10310
rect 10670 10308 10694 10310
rect 10750 10308 10774 10310
rect 10830 10308 10854 10310
rect 10910 10308 10916 10310
rect 10608 10299 10916 10308
rect 11164 9586 11192 10610
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 9994 11284 10406
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11268 9820 11576 9829
rect 11268 9818 11274 9820
rect 11330 9818 11354 9820
rect 11410 9818 11434 9820
rect 11490 9818 11514 9820
rect 11570 9818 11576 9820
rect 11330 9766 11332 9818
rect 11512 9766 11514 9818
rect 11268 9764 11274 9766
rect 11330 9764 11354 9766
rect 11410 9764 11434 9766
rect 11490 9764 11514 9766
rect 11570 9764 11576 9766
rect 11268 9755 11576 9764
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10608 9276 10916 9285
rect 10608 9274 10614 9276
rect 10670 9274 10694 9276
rect 10750 9274 10774 9276
rect 10830 9274 10854 9276
rect 10910 9274 10916 9276
rect 10670 9222 10672 9274
rect 10852 9222 10854 9274
rect 10608 9220 10614 9222
rect 10670 9220 10694 9222
rect 10750 9220 10774 9222
rect 10830 9220 10854 9222
rect 10910 9220 10916 9222
rect 10608 9211 10916 9220
rect 11058 9208 11114 9217
rect 11058 9143 11060 9152
rect 11112 9143 11114 9152
rect 11060 9114 11112 9120
rect 10782 8936 10838 8945
rect 10782 8871 10784 8880
rect 10836 8871 10838 8880
rect 10784 8842 10836 8848
rect 11268 8732 11576 8741
rect 11268 8730 11274 8732
rect 11330 8730 11354 8732
rect 11410 8730 11434 8732
rect 11490 8730 11514 8732
rect 11570 8730 11576 8732
rect 11330 8678 11332 8730
rect 11512 8678 11514 8730
rect 11268 8676 11274 8678
rect 11330 8676 11354 8678
rect 11410 8676 11434 8678
rect 11490 8676 11514 8678
rect 11570 8676 11576 8678
rect 11268 8667 11576 8676
rect 10608 8188 10916 8197
rect 10608 8186 10614 8188
rect 10670 8186 10694 8188
rect 10750 8186 10774 8188
rect 10830 8186 10854 8188
rect 10910 8186 10916 8188
rect 10670 8134 10672 8186
rect 10852 8134 10854 8186
rect 10608 8132 10614 8134
rect 10670 8132 10694 8134
rect 10750 8132 10774 8134
rect 10830 8132 10854 8134
rect 10910 8132 10916 8134
rect 10608 8123 10916 8132
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10704 7342 10732 7754
rect 10600 7336 10652 7342
rect 10598 7304 10600 7313
rect 10692 7336 10744 7342
rect 10652 7304 10654 7313
rect 10692 7278 10744 7284
rect 10598 7239 10654 7248
rect 10608 7100 10916 7109
rect 10608 7098 10614 7100
rect 10670 7098 10694 7100
rect 10750 7098 10774 7100
rect 10830 7098 10854 7100
rect 10910 7098 10916 7100
rect 10670 7046 10672 7098
rect 10852 7046 10854 7098
rect 10608 7044 10614 7046
rect 10670 7044 10694 7046
rect 10750 7044 10774 7046
rect 10830 7044 10854 7046
rect 10910 7044 10916 7046
rect 10608 7035 10916 7044
rect 10980 6934 11008 7958
rect 11624 7834 11652 12406
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11218 11836 12174
rect 12084 11218 12112 12854
rect 12268 12850 12296 14282
rect 12820 14278 12848 16934
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13530 12848 14214
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12530 13424 12586 13433
rect 12530 13359 12532 13368
rect 12584 13359 12586 13368
rect 12532 13330 12584 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12360 12238 12388 13262
rect 12808 12436 12860 12442
rect 12912 12434 12940 16526
rect 13084 16176 13136 16182
rect 13188 16153 13216 17167
rect 13556 17082 13584 17614
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13556 17066 13676 17082
rect 13556 17060 13688 17066
rect 13556 17054 13636 17060
rect 13556 16794 13584 17054
rect 13636 17002 13688 17008
rect 13740 16998 13768 17138
rect 14016 16998 14044 17614
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13084 16118 13136 16124
rect 13174 16144 13230 16153
rect 13096 15706 13124 16118
rect 13174 16079 13230 16088
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 15502 13216 16079
rect 13176 15496 13228 15502
rect 13228 15456 13308 15484
rect 13176 15438 13228 15444
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 12889 13124 14962
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13082 12880 13138 12889
rect 13188 12850 13216 13738
rect 13280 13326 13308 15456
rect 13636 14408 13688 14414
rect 13740 14396 13768 16934
rect 14108 16658 14136 17206
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 16250 14136 16594
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15570 13952 15846
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13688 14368 13768 14396
rect 13636 14350 13688 14356
rect 13648 14074 13676 14350
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 14074 14136 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13556 13530 13584 13942
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13082 12815 13138 12824
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13280 12714 13308 12922
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13464 12646 13492 12854
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 12860 12406 12940 12434
rect 14200 12434 14228 18158
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16250 14320 16390
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14384 14822 14412 17614
rect 14752 16590 14780 20946
rect 15304 20942 15332 21490
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14936 18834 14964 19722
rect 15120 18873 15148 20810
rect 15304 19334 15332 20878
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15212 19306 15332 19334
rect 15106 18864 15162 18873
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 15028 18822 15106 18850
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14844 17338 14872 18158
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14832 16448 14884 16454
rect 14660 16408 14832 16436
rect 14660 16250 14688 16408
rect 14884 16408 14964 16436
rect 14832 16390 14884 16396
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14752 14822 14780 15438
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14200 12406 14320 12434
rect 12808 12378 12860 12384
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11218 12388 11494
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 11808 10674 11836 11154
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10810 13124 11018
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11716 8906 11744 10542
rect 12084 10266 12112 10542
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 13648 10062 13676 10950
rect 13740 10198 13768 11630
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 11900 9382 11928 9930
rect 12452 9654 12480 9930
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9110 12848 9318
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12912 8906 12940 9862
rect 12990 9208 13046 9217
rect 13084 9172 13136 9178
rect 13046 9152 13084 9160
rect 12990 9143 13084 9152
rect 13004 9132 13084 9143
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11164 7806 11652 7834
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11704 7812 11756 7818
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10612 6458 10640 6870
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6458 10732 6734
rect 11072 6730 11100 7754
rect 11164 7290 11192 7806
rect 11704 7754 11756 7760
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11268 7644 11576 7653
rect 11268 7642 11274 7644
rect 11330 7642 11354 7644
rect 11410 7642 11434 7644
rect 11490 7642 11514 7644
rect 11570 7642 11576 7644
rect 11330 7590 11332 7642
rect 11512 7590 11514 7642
rect 11268 7588 11274 7590
rect 11330 7588 11354 7590
rect 11410 7588 11434 7590
rect 11490 7588 11514 7590
rect 11570 7588 11576 7590
rect 11268 7579 11576 7588
rect 11164 7262 11284 7290
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11256 6746 11284 7262
rect 11624 6866 11652 7686
rect 11716 7002 11744 7754
rect 11900 7546 11928 7822
rect 11992 7546 12020 8026
rect 12084 7886 12112 8774
rect 12820 8566 12848 8774
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11794 7440 11850 7449
rect 11794 7375 11796 7384
rect 11848 7375 11850 7384
rect 11796 7346 11848 7352
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11808 6934 11836 7346
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11164 6718 11284 6746
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10608 6012 10916 6021
rect 10608 6010 10614 6012
rect 10670 6010 10694 6012
rect 10750 6010 10774 6012
rect 10830 6010 10854 6012
rect 10910 6010 10916 6012
rect 10670 5958 10672 6010
rect 10852 5958 10854 6010
rect 10608 5956 10614 5958
rect 10670 5956 10694 5958
rect 10750 5956 10774 5958
rect 10830 5956 10854 5958
rect 10910 5956 10916 5958
rect 10608 5947 10916 5956
rect 10152 5766 10548 5794
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6380 3058 6408 3334
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 4169 2748 4477 2757
rect 4169 2746 4175 2748
rect 4231 2746 4255 2748
rect 4311 2746 4335 2748
rect 4391 2746 4415 2748
rect 4471 2746 4477 2748
rect 4231 2694 4233 2746
rect 4413 2694 4415 2746
rect 4169 2692 4175 2694
rect 4231 2692 4255 2694
rect 4311 2692 4335 2694
rect 4391 2692 4415 2694
rect 4471 2692 4477 2694
rect 4169 2683 4477 2692
rect 5552 2650 5580 2858
rect 6564 2854 6592 4082
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3058 6684 3946
rect 6748 3942 6776 4082
rect 8036 4078 8064 4558
rect 8312 4214 8340 4626
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5736 2446 5764 2790
rect 6748 2774 6776 3878
rect 8312 3602 8340 4150
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 6932 3194 6960 3402
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7392 3058 7420 3334
rect 8036 3194 8064 3402
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 8312 2990 8340 3538
rect 8404 3534 8432 4558
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8404 3074 8432 3470
rect 8496 3194 8524 4014
rect 8864 3194 8892 4150
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3534 9628 3946
rect 9784 3942 9812 4014
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3534 9812 3878
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9140 3126 9168 3334
rect 9128 3120 9180 3126
rect 8404 3058 8708 3074
rect 9128 3062 9180 3068
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 8392 3052 8720 3058
rect 8444 3046 8668 3052
rect 8392 2994 8444 3000
rect 8668 2994 8720 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 6656 2746 6776 2774
rect 6656 2446 6684 2746
rect 8956 2446 8984 2994
rect 9784 2650 9812 3062
rect 9968 2990 9996 4422
rect 10060 4282 10088 4558
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10152 2514 10180 5766
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4690 10548 4966
rect 10608 4924 10916 4933
rect 10608 4922 10614 4924
rect 10670 4922 10694 4924
rect 10750 4922 10774 4924
rect 10830 4922 10854 4924
rect 10910 4922 10916 4924
rect 10670 4870 10672 4922
rect 10852 4870 10854 4922
rect 10608 4868 10614 4870
rect 10670 4868 10694 4870
rect 10750 4868 10774 4870
rect 10830 4868 10854 4870
rect 10910 4868 10916 4870
rect 10608 4859 10916 4868
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 3738 10272 4422
rect 10416 4140 10468 4146
rect 10520 4128 10548 4626
rect 11072 4593 11100 4762
rect 11058 4584 11114 4593
rect 11058 4519 11114 4528
rect 10468 4100 10548 4128
rect 10416 4082 10468 4088
rect 11072 4078 11100 4519
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10428 3602 10456 3878
rect 10608 3836 10916 3845
rect 10608 3834 10614 3836
rect 10670 3834 10694 3836
rect 10750 3834 10774 3836
rect 10830 3834 10854 3836
rect 10910 3834 10916 3836
rect 10670 3782 10672 3834
rect 10852 3782 10854 3834
rect 10608 3780 10614 3782
rect 10670 3780 10694 3782
rect 10750 3780 10774 3782
rect 10830 3780 10854 3782
rect 10910 3780 10916 3782
rect 10608 3771 10916 3780
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 11072 3194 11100 4014
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10608 2748 10916 2757
rect 10608 2746 10614 2748
rect 10670 2746 10694 2748
rect 10750 2746 10774 2748
rect 10830 2746 10854 2748
rect 10910 2746 10916 2748
rect 10670 2694 10672 2746
rect 10852 2694 10854 2746
rect 10608 2692 10614 2694
rect 10670 2692 10694 2694
rect 10750 2692 10774 2694
rect 10830 2692 10854 2694
rect 10910 2692 10916 2694
rect 10608 2683 10916 2692
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 11164 2446 11192 6718
rect 11992 6662 12020 6938
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11268 6556 11576 6565
rect 11268 6554 11274 6556
rect 11330 6554 11354 6556
rect 11410 6554 11434 6556
rect 11490 6554 11514 6556
rect 11570 6554 11576 6556
rect 11330 6502 11332 6554
rect 11512 6502 11514 6554
rect 11268 6500 11274 6502
rect 11330 6500 11354 6502
rect 11410 6500 11434 6502
rect 11490 6500 11514 6502
rect 11570 6500 11576 6502
rect 11268 6491 11576 6500
rect 11268 5468 11576 5477
rect 11268 5466 11274 5468
rect 11330 5466 11354 5468
rect 11410 5466 11434 5468
rect 11490 5466 11514 5468
rect 11570 5466 11576 5468
rect 11330 5414 11332 5466
rect 11512 5414 11514 5466
rect 11268 5412 11274 5414
rect 11330 5412 11354 5414
rect 11410 5412 11434 5414
rect 11490 5412 11514 5414
rect 11570 5412 11576 5414
rect 11268 5403 11576 5412
rect 12176 5098 12204 7142
rect 12452 6798 12480 7686
rect 12728 7546 12756 7958
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12912 5914 12940 8298
rect 13004 8090 13032 9132
rect 13084 9114 13136 9120
rect 13648 9110 13676 9998
rect 13740 9178 13768 10134
rect 14200 10062 14228 10950
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13266 8936 13322 8945
rect 13176 8900 13228 8906
rect 13322 8880 13492 8888
rect 13266 8871 13268 8880
rect 13176 8842 13228 8848
rect 13320 8860 13492 8880
rect 13268 8842 13320 8848
rect 13188 8634 13216 8842
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13464 8566 13492 8860
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13004 7274 13032 8026
rect 13096 7886 13124 8434
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8090 13400 8230
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7954 13492 8502
rect 13648 8498 13676 9046
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13648 8090 13676 8434
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 13096 6798 13124 7822
rect 13464 7478 13492 7890
rect 13648 7886 13676 8026
rect 13740 7954 13768 8570
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13648 7410 13676 7822
rect 13740 7546 13768 7890
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13004 5914 13032 6666
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13372 5642 13400 6598
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13464 5234 13492 7142
rect 13556 6934 13584 7142
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13832 6798 13860 9318
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14108 8430 14136 9114
rect 14200 8634 14228 9998
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14096 8424 14148 8430
rect 14016 8384 14096 8412
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13924 5846 13952 8230
rect 14016 7478 14044 8384
rect 14096 8366 14148 8372
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 8090 14136 8230
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14200 7274 14228 7482
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13636 5296 13688 5302
rect 13634 5264 13636 5273
rect 13688 5264 13690 5273
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13452 5228 13504 5234
rect 13634 5199 13690 5208
rect 13452 5170 13504 5176
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 11268 4380 11576 4389
rect 11268 4378 11274 4380
rect 11330 4378 11354 4380
rect 11410 4378 11434 4380
rect 11490 4378 11514 4380
rect 11570 4378 11576 4380
rect 11330 4326 11332 4378
rect 11512 4326 11514 4378
rect 11268 4324 11274 4326
rect 11330 4324 11354 4326
rect 11410 4324 11434 4326
rect 11490 4324 11514 4326
rect 11570 4324 11576 4326
rect 11268 4315 11576 4324
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3466 11652 3878
rect 12176 3738 12204 5034
rect 12452 4146 12480 5170
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4282 12572 4422
rect 12636 4282 12664 5170
rect 13096 5030 13124 5170
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4758 13124 4966
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13096 4622 13124 4694
rect 13280 4622 13308 5034
rect 13464 4808 13492 5170
rect 13924 5166 13952 5782
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13544 4820 13596 4826
rect 13464 4780 13544 4808
rect 13544 4762 13596 4768
rect 13084 4616 13136 4622
rect 13082 4584 13084 4593
rect 13268 4616 13320 4622
rect 13136 4584 13138 4593
rect 12900 4548 12952 4554
rect 13268 4558 13320 4564
rect 13082 4519 13138 4528
rect 12900 4490 12952 4496
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12544 3466 12572 4218
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12728 3534 12756 4082
rect 12912 4078 12940 4490
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4214 13032 4422
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 13360 4208 13412 4214
rect 13556 4196 13584 4762
rect 13924 4622 13952 5102
rect 14016 5030 14044 5170
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 4282 13952 4422
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14108 4214 14136 4558
rect 13412 4168 13584 4196
rect 13360 4150 13412 4156
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13004 3602 13032 4150
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13372 3534 13400 3878
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13464 3466 13492 3946
rect 13556 3738 13584 4168
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 14108 3398 14136 4150
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 11268 3292 11576 3301
rect 11268 3290 11274 3292
rect 11330 3290 11354 3292
rect 11410 3290 11434 3292
rect 11490 3290 11514 3292
rect 11570 3290 11576 3292
rect 11330 3238 11332 3290
rect 11512 3238 11514 3290
rect 11268 3236 11274 3238
rect 11330 3236 11354 3238
rect 11410 3236 11434 3238
rect 11490 3236 11514 3238
rect 11570 3236 11576 3238
rect 11268 3227 11576 3236
rect 14292 2446 14320 12406
rect 14384 6905 14412 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14074 14596 14418
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14462 12744 14518 12753
rect 14462 12679 14518 12688
rect 14476 12434 14504 12679
rect 14476 12406 14596 12434
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14476 10742 14504 11834
rect 14568 11694 14596 12406
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 10198 14504 10542
rect 14568 10266 14596 11086
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14476 8566 14504 10134
rect 14660 9586 14688 12174
rect 14752 10606 14780 14758
rect 14936 14414 14964 16408
rect 15028 16130 15056 18822
rect 15106 18799 15162 18808
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15120 18426 15148 18702
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15212 16810 15240 19306
rect 15396 18970 15424 20334
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15488 18766 15516 19178
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15304 17270 15332 18702
rect 15488 18086 15516 18702
rect 15580 18630 15608 19790
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18426 15608 18566
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15474 17912 15530 17921
rect 15474 17847 15476 17856
rect 15528 17847 15530 17856
rect 15476 17818 15528 17824
rect 15672 17678 15700 20810
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15842 20360 15898 20369
rect 15842 20295 15898 20304
rect 15856 19854 15884 20295
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15764 18766 15792 19790
rect 15948 19242 15976 20402
rect 16488 20392 16540 20398
rect 16394 20360 16450 20369
rect 16488 20334 16540 20340
rect 16394 20295 16396 20304
rect 16448 20295 16450 20304
rect 16396 20266 16448 20272
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 20058 16160 20198
rect 16500 20058 16528 20334
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15752 18760 15804 18766
rect 15804 18708 15884 18714
rect 15752 18702 15884 18708
rect 15764 18686 15884 18702
rect 15948 18698 15976 18838
rect 15856 18290 15884 18686
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18442 15976 18634
rect 16040 18630 16068 19654
rect 16224 18970 16252 19790
rect 16408 19242 16436 19790
rect 16592 19530 16620 22086
rect 16684 19922 16712 22578
rect 16764 22432 16816 22438
rect 16816 22380 16896 22386
rect 16764 22374 16896 22380
rect 16776 22358 16896 22374
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16776 22030 16804 22170
rect 16868 22098 16896 22358
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16500 19514 16620 19530
rect 16488 19508 16620 19514
rect 16540 19502 16620 19508
rect 16488 19450 16540 19456
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16408 18766 16436 19178
rect 16500 18902 16528 19314
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 15948 18414 16068 18442
rect 16224 18426 16252 18566
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15764 17814 15792 18226
rect 15948 18170 15976 18226
rect 15856 18142 15976 18170
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15382 17368 15438 17377
rect 15382 17303 15384 17312
rect 15436 17303 15438 17312
rect 15384 17274 15436 17280
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15212 16782 15332 16810
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15028 16102 15148 16130
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15706 15056 15982
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15120 14618 15148 16102
rect 15212 15706 15240 16662
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14924 14408 14976 14414
rect 14976 14368 15056 14396
rect 14924 14350 14976 14356
rect 14844 13734 14872 14350
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 14074 14964 14214
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15028 14006 15056 14368
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13326 14872 13670
rect 14936 13326 14964 13874
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13530 15056 13806
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14924 13320 14976 13326
rect 15304 13274 15332 16782
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13530 15424 13670
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 14924 13262 14976 13268
rect 15212 13246 15332 13274
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12782 15056 13126
rect 15016 12776 15068 12782
rect 15108 12776 15160 12782
rect 15016 12718 15068 12724
rect 15106 12744 15108 12753
rect 15160 12744 15162 12753
rect 15106 12679 15162 12688
rect 15212 11801 15240 13246
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12850 15332 13126
rect 15488 12918 15516 15438
rect 15672 14385 15700 17070
rect 15856 17066 15884 18142
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 16794 15792 16934
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15658 14376 15714 14385
rect 15658 14311 15660 14320
rect 15712 14311 15714 14320
rect 15660 14282 15712 14288
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15580 12986 15608 14214
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12986 15792 13194
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 11898 15332 12786
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 12306 15424 12582
rect 15764 12306 15792 12650
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 15212 10606 15240 11727
rect 15396 11200 15424 12242
rect 15568 11212 15620 11218
rect 15396 11172 15568 11200
rect 15568 11154 15620 11160
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15672 10810 15700 11018
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10062 15240 10542
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 8634 15056 9454
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14464 8560 14516 8566
rect 14516 8520 14596 8548
rect 14464 8502 14516 8508
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 7342 14504 7754
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14568 7274 14596 8520
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7546 14688 7822
rect 14844 7818 14872 8230
rect 15028 7886 15056 8298
rect 15120 7886 15148 8774
rect 15304 8498 15332 10610
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15580 9178 15608 9590
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15396 8430 15424 8842
rect 15764 8566 15792 9318
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14370 6896 14426 6905
rect 14370 6831 14426 6840
rect 14384 5574 14412 6831
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14384 4457 14412 4490
rect 14370 4448 14426 4457
rect 14370 4383 14426 4392
rect 14384 3466 14412 4383
rect 14752 3942 14780 7754
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15120 7206 15148 7686
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15212 6769 15240 7686
rect 15198 6760 15254 6769
rect 15198 6695 15254 6704
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5642 15056 6054
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15106 5264 15162 5273
rect 15106 5199 15108 5208
rect 15160 5199 15162 5208
rect 15108 5170 15160 5176
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15028 4622 15056 4966
rect 15120 4690 15148 4966
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14936 4078 14964 4558
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3194 14872 3402
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15212 3058 15240 6258
rect 15396 6254 15424 8366
rect 15764 7886 15792 8502
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15488 4214 15516 7754
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 4826 15608 5646
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15488 3942 15516 4150
rect 15672 4146 15700 4422
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15856 2446 15884 17002
rect 15948 15314 15976 18022
rect 16040 17898 16068 18414
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16408 18086 16436 18702
rect 16592 18154 16620 19382
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16040 17870 16436 17898
rect 16684 17882 16712 19858
rect 16776 19446 16804 21558
rect 16960 21146 16988 22714
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17047 22332 17355 22341
rect 17047 22330 17053 22332
rect 17109 22330 17133 22332
rect 17189 22330 17213 22332
rect 17269 22330 17293 22332
rect 17349 22330 17355 22332
rect 17109 22278 17111 22330
rect 17291 22278 17293 22330
rect 17047 22276 17053 22278
rect 17109 22276 17133 22278
rect 17189 22276 17213 22278
rect 17269 22276 17293 22278
rect 17349 22276 17355 22278
rect 17047 22267 17355 22276
rect 17972 22098 18000 22646
rect 18050 22128 18106 22137
rect 17960 22092 18012 22098
rect 18050 22063 18106 22072
rect 17960 22034 18012 22040
rect 18064 22030 18092 22063
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17604 21486 17632 21966
rect 17707 21788 18015 21797
rect 17707 21786 17713 21788
rect 17769 21786 17793 21788
rect 17849 21786 17873 21788
rect 17929 21786 17953 21788
rect 18009 21786 18015 21788
rect 17769 21734 17771 21786
rect 17951 21734 17953 21786
rect 17707 21732 17713 21734
rect 17769 21732 17793 21734
rect 17849 21732 17873 21734
rect 17929 21732 17953 21734
rect 18009 21732 18015 21734
rect 17707 21723 18015 21732
rect 18064 21554 18092 21966
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18248 21554 18276 21830
rect 18340 21690 18368 23054
rect 18524 22234 18552 23054
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18616 21962 18644 22510
rect 18800 22094 18828 22510
rect 19076 22234 19104 23054
rect 19628 22982 19656 23820
rect 19800 23802 19852 23808
rect 19904 23730 19932 24822
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24342 20116 24754
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19904 23322 19932 23666
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19720 23118 19748 23258
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19892 23044 19944 23050
rect 19892 22986 19944 22992
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 19812 22574 19840 22918
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19720 22420 19748 22510
rect 19904 22420 19932 22986
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19720 22392 19932 22420
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18708 22066 18828 22094
rect 18708 22030 18736 22066
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18708 21894 18736 21966
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17047 21244 17355 21253
rect 17047 21242 17053 21244
rect 17109 21242 17133 21244
rect 17189 21242 17213 21244
rect 17269 21242 17293 21244
rect 17349 21242 17355 21244
rect 17109 21190 17111 21242
rect 17291 21190 17293 21242
rect 17047 21188 17053 21190
rect 17109 21188 17133 21190
rect 17189 21188 17213 21190
rect 17269 21188 17293 21190
rect 17349 21188 17355 21190
rect 17047 21179 17355 21188
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17052 20505 17080 20538
rect 17420 20534 17448 20742
rect 17408 20528 17460 20534
rect 17038 20496 17094 20505
rect 16856 20460 16908 20466
rect 17408 20470 17460 20476
rect 17038 20431 17040 20440
rect 16856 20402 16908 20408
rect 17092 20431 17094 20440
rect 17040 20402 17092 20408
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16868 19394 16896 20402
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16960 19514 16988 20266
rect 17047 20156 17355 20165
rect 17047 20154 17053 20156
rect 17109 20154 17133 20156
rect 17189 20154 17213 20156
rect 17269 20154 17293 20156
rect 17349 20154 17355 20156
rect 17109 20102 17111 20154
rect 17291 20102 17293 20154
rect 17047 20100 17053 20102
rect 17109 20100 17133 20102
rect 17189 20100 17213 20102
rect 17269 20100 17293 20102
rect 17349 20100 17355 20102
rect 17047 20091 17355 20100
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17052 19394 17080 19790
rect 16868 19366 17080 19394
rect 16764 19304 16816 19310
rect 16868 19258 16896 19366
rect 16816 19252 16896 19258
rect 16764 19246 16896 19252
rect 16776 19230 16896 19246
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16776 18902 16804 19110
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16868 18766 16896 19110
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16868 18290 16896 18702
rect 16960 18426 16988 19366
rect 17047 19068 17355 19077
rect 17047 19066 17053 19068
rect 17109 19066 17133 19068
rect 17189 19066 17213 19068
rect 17269 19066 17293 19068
rect 17349 19066 17355 19068
rect 17109 19014 17111 19066
rect 17291 19014 17293 19066
rect 17047 19012 17053 19014
rect 17109 19012 17133 19014
rect 17189 19012 17213 19014
rect 17269 19012 17293 19014
rect 17349 19012 17355 19014
rect 17047 19003 17355 19012
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 17052 18170 17080 18566
rect 17328 18426 17356 18906
rect 17420 18698 17448 20470
rect 17512 20398 17540 20878
rect 17604 20482 17632 21422
rect 18800 21350 18828 21966
rect 18984 21622 19012 22170
rect 19904 22098 19932 22392
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19996 21894 20024 22646
rect 20088 22234 20116 23258
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20180 22094 20208 25842
rect 21284 24886 21312 26250
rect 24146 26140 24454 26149
rect 24146 26138 24152 26140
rect 24208 26138 24232 26140
rect 24288 26138 24312 26140
rect 24368 26138 24392 26140
rect 24448 26138 24454 26140
rect 24208 26086 24210 26138
rect 24390 26086 24392 26138
rect 24146 26084 24152 26086
rect 24208 26084 24232 26086
rect 24288 26084 24312 26086
rect 24368 26084 24392 26086
rect 24448 26084 24454 26086
rect 24146 26075 24454 26084
rect 23486 25596 23794 25605
rect 23486 25594 23492 25596
rect 23548 25594 23572 25596
rect 23628 25594 23652 25596
rect 23708 25594 23732 25596
rect 23788 25594 23794 25596
rect 23548 25542 23550 25594
rect 23730 25542 23732 25594
rect 23486 25540 23492 25542
rect 23548 25540 23572 25542
rect 23628 25540 23652 25542
rect 23708 25540 23732 25542
rect 23788 25540 23794 25542
rect 23486 25531 23794 25540
rect 24146 25052 24454 25061
rect 24146 25050 24152 25052
rect 24208 25050 24232 25052
rect 24288 25050 24312 25052
rect 24368 25050 24392 25052
rect 24448 25050 24454 25052
rect 24208 24998 24210 25050
rect 24390 24998 24392 25050
rect 24146 24996 24152 24998
rect 24208 24996 24232 24998
rect 24288 24996 24312 24998
rect 24368 24996 24392 24998
rect 24448 24996 24454 24998
rect 24146 24987 24454 24996
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20456 23118 20484 24210
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23662 20668 24074
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 21284 23712 21312 24142
rect 21456 23724 21508 23730
rect 21284 23684 21456 23712
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20916 23322 20944 23666
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 21284 23050 21312 23684
rect 21456 23666 21508 23672
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 20548 22506 20576 22986
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20548 22234 20576 22442
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20088 22066 20208 22094
rect 20088 22030 20116 22066
rect 20640 22030 20668 22578
rect 20732 22438 20760 22986
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20824 22642 20852 22918
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20824 22098 20852 22578
rect 21376 22234 21404 23054
rect 21560 22574 21588 23666
rect 21652 23118 21680 24686
rect 22204 24342 22232 24686
rect 22572 24410 22600 24822
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21928 23798 21956 24006
rect 22204 23866 22232 24278
rect 23308 24274 23336 24550
rect 23486 24508 23794 24517
rect 23486 24506 23492 24508
rect 23548 24506 23572 24508
rect 23628 24506 23652 24508
rect 23708 24506 23732 24508
rect 23788 24506 23794 24508
rect 23548 24454 23550 24506
rect 23730 24454 23732 24506
rect 23486 24452 23492 24454
rect 23548 24452 23572 24454
rect 23628 24452 23652 24454
rect 23708 24452 23732 24454
rect 23788 24452 23794 24454
rect 23486 24443 23794 24452
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 22664 23730 22692 24142
rect 24146 23964 24454 23973
rect 24146 23962 24152 23964
rect 24208 23962 24232 23964
rect 24288 23962 24312 23964
rect 24368 23962 24392 23964
rect 24448 23962 24454 23964
rect 24208 23910 24210 23962
rect 24390 23910 24392 23962
rect 24146 23908 24152 23910
rect 24208 23908 24232 23910
rect 24288 23908 24312 23910
rect 24368 23908 24392 23910
rect 24448 23908 24454 23910
rect 24146 23899 24454 23908
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22664 23610 22692 23666
rect 22572 23582 22692 23610
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22112 23322 22140 23462
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22296 23186 22324 23462
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22710 21680 23054
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22710 22140 22918
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21560 22098 21588 22374
rect 21652 22166 21680 22510
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21652 22030 21680 22102
rect 22572 22030 22600 23582
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22664 23050 22692 23462
rect 23486 23420 23794 23429
rect 23486 23418 23492 23420
rect 23548 23418 23572 23420
rect 23628 23418 23652 23420
rect 23708 23418 23732 23420
rect 23788 23418 23794 23420
rect 23548 23366 23550 23418
rect 23730 23366 23732 23418
rect 23486 23364 23492 23366
rect 23548 23364 23572 23366
rect 23628 23364 23652 23366
rect 23708 23364 23732 23366
rect 23788 23364 23794 23366
rect 23486 23355 23794 23364
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 24146 22876 24454 22885
rect 24146 22874 24152 22876
rect 24208 22874 24232 22876
rect 24288 22874 24312 22876
rect 24368 22874 24392 22876
rect 24448 22874 24454 22876
rect 24208 22822 24210 22874
rect 24390 22822 24392 22874
rect 24146 22820 24152 22822
rect 24208 22820 24232 22822
rect 24288 22820 24312 22822
rect 24368 22820 24392 22822
rect 24448 22820 24454 22822
rect 24146 22811 24454 22820
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22664 22098 22692 22646
rect 23486 22332 23794 22341
rect 23486 22330 23492 22332
rect 23548 22330 23572 22332
rect 23628 22330 23652 22332
rect 23708 22330 23732 22332
rect 23788 22330 23794 22332
rect 23548 22278 23550 22330
rect 23730 22278 23732 22330
rect 23486 22276 23492 22278
rect 23548 22276 23572 22278
rect 23628 22276 23652 22278
rect 23708 22276 23732 22278
rect 23788 22276 23794 22278
rect 23486 22267 23794 22276
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 20088 21894 20116 21966
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 20088 21486 20116 21830
rect 24146 21788 24454 21797
rect 24146 21786 24152 21788
rect 24208 21786 24232 21788
rect 24288 21786 24312 21788
rect 24368 21786 24392 21788
rect 24448 21786 24454 21788
rect 24208 21734 24210 21786
rect 24390 21734 24392 21786
rect 24146 21732 24152 21734
rect 24208 21732 24232 21734
rect 24288 21732 24312 21734
rect 24368 21732 24392 21734
rect 24448 21732 24454 21734
rect 24146 21723 24454 21732
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 23486 21244 23794 21253
rect 23486 21242 23492 21244
rect 23548 21242 23572 21244
rect 23628 21242 23652 21244
rect 23708 21242 23732 21244
rect 23788 21242 23794 21244
rect 23548 21190 23550 21242
rect 23730 21190 23732 21242
rect 23486 21188 23492 21190
rect 23548 21188 23572 21190
rect 23628 21188 23652 21190
rect 23708 21188 23732 21190
rect 23788 21188 23794 21190
rect 23486 21179 23794 21188
rect 17707 20700 18015 20709
rect 17707 20698 17713 20700
rect 17769 20698 17793 20700
rect 17849 20698 17873 20700
rect 17929 20698 17953 20700
rect 18009 20698 18015 20700
rect 17769 20646 17771 20698
rect 17951 20646 17953 20698
rect 17707 20644 17713 20646
rect 17769 20644 17793 20646
rect 17849 20644 17873 20646
rect 17929 20644 17953 20646
rect 18009 20644 18015 20646
rect 17707 20635 18015 20644
rect 24146 20700 24454 20709
rect 24146 20698 24152 20700
rect 24208 20698 24232 20700
rect 24288 20698 24312 20700
rect 24368 20698 24392 20700
rect 24448 20698 24454 20700
rect 24208 20646 24210 20698
rect 24390 20646 24392 20698
rect 24146 20644 24152 20646
rect 24208 20644 24232 20646
rect 24288 20644 24312 20646
rect 24368 20644 24392 20646
rect 24448 20644 24454 20646
rect 24146 20635 24454 20644
rect 24596 20602 24624 27338
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 18604 20528 18656 20534
rect 17604 20454 17816 20482
rect 18604 20470 18656 20476
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17512 20074 17540 20334
rect 17512 20046 17632 20074
rect 17696 20058 17724 20334
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 16868 18142 17080 18170
rect 16868 18086 16896 18142
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 15502 16344 16390
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 15948 15286 16344 15314
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 13190 15976 14554
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13394 16160 14214
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15948 12918 15976 13126
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 16132 12850 16160 13126
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12434 16252 12582
rect 16132 12406 16252 12434
rect 16132 11830 16160 12406
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 15948 11354 15976 11766
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16040 11150 16068 11222
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 8974 16068 11086
rect 16316 9674 16344 15286
rect 16224 9646 16344 9674
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16224 6304 16252 9646
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 6458 16344 6734
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16224 6276 16344 6304
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16224 4214 16252 4558
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16118 4040 16174 4049
rect 16118 3975 16120 3984
rect 16172 3975 16174 3984
rect 16120 3946 16172 3952
rect 16224 3738 16252 4150
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16316 2514 16344 6276
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16408 2378 16436 17870
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 16266 16620 16594
rect 16500 16238 16620 16266
rect 16500 15434 16528 16238
rect 16684 16182 16712 16934
rect 16776 16590 16804 17138
rect 16960 16674 16988 18022
rect 17047 17980 17355 17989
rect 17047 17978 17053 17980
rect 17109 17978 17133 17980
rect 17189 17978 17213 17980
rect 17269 17978 17293 17980
rect 17349 17978 17355 17980
rect 17109 17926 17111 17978
rect 17291 17926 17293 17978
rect 17047 17924 17053 17926
rect 17109 17924 17133 17926
rect 17189 17924 17213 17926
rect 17269 17924 17293 17926
rect 17349 17924 17355 17926
rect 17047 17915 17355 17924
rect 17047 16892 17355 16901
rect 17047 16890 17053 16892
rect 17109 16890 17133 16892
rect 17189 16890 17213 16892
rect 17269 16890 17293 16892
rect 17349 16890 17355 16892
rect 17109 16838 17111 16890
rect 17291 16838 17293 16890
rect 17047 16836 17053 16838
rect 17109 16836 17133 16838
rect 17189 16836 17213 16838
rect 17269 16836 17293 16838
rect 17349 16836 17355 16838
rect 17047 16827 17355 16836
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 16868 16646 16988 16674
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16868 16522 16896 16646
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16960 16182 16988 16458
rect 17052 16182 17080 16730
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 17040 16176 17092 16182
rect 17420 16153 17448 16526
rect 17040 16118 17092 16124
rect 17406 16144 17462 16153
rect 16580 16108 16632 16114
rect 17406 16079 17462 16088
rect 16580 16050 16632 16056
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16592 15162 16620 16050
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16684 15162 16712 15370
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16592 14618 16620 15098
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16580 14408 16632 14414
rect 16684 14396 16712 15098
rect 16776 15094 16804 15982
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16868 15638 16896 15846
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16868 15026 16896 15574
rect 16960 15570 16988 15846
rect 17047 15804 17355 15813
rect 17047 15802 17053 15804
rect 17109 15802 17133 15804
rect 17189 15802 17213 15804
rect 17269 15802 17293 15804
rect 17349 15802 17355 15804
rect 17109 15750 17111 15802
rect 17291 15750 17293 15802
rect 17047 15748 17053 15750
rect 17109 15748 17133 15750
rect 17189 15748 17213 15750
rect 17269 15748 17293 15750
rect 17349 15748 17355 15750
rect 17047 15739 17355 15748
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16868 14414 16896 14962
rect 16632 14368 16712 14396
rect 16856 14408 16908 14414
rect 16580 14350 16632 14356
rect 16856 14350 16908 14356
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16500 11218 16528 11630
rect 16684 11558 16712 14214
rect 16960 13734 16988 15030
rect 17047 14716 17355 14725
rect 17047 14714 17053 14716
rect 17109 14714 17133 14716
rect 17189 14714 17213 14716
rect 17269 14714 17293 14716
rect 17349 14714 17355 14716
rect 17109 14662 17111 14714
rect 17291 14662 17293 14714
rect 17047 14660 17053 14662
rect 17109 14660 17133 14662
rect 17189 14660 17213 14662
rect 17269 14660 17293 14662
rect 17349 14660 17355 14662
rect 17047 14651 17355 14660
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17236 14521 17264 14554
rect 17222 14512 17278 14521
rect 17222 14447 17278 14456
rect 17420 14414 17448 15914
rect 17512 15706 17540 19858
rect 17604 19854 17632 20046
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17788 19938 17816 20454
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18432 20058 18460 20334
rect 18616 20058 18644 20470
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 17788 19910 18276 19938
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17604 18850 17632 19790
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17707 19612 18015 19621
rect 17707 19610 17713 19612
rect 17769 19610 17793 19612
rect 17849 19610 17873 19612
rect 17929 19610 17953 19612
rect 18009 19610 18015 19612
rect 17769 19558 17771 19610
rect 17951 19558 17953 19610
rect 17707 19556 17713 19558
rect 17769 19556 17793 19558
rect 17849 19556 17873 19558
rect 17929 19556 17953 19558
rect 18009 19556 18015 19558
rect 17707 19547 18015 19556
rect 18064 19310 18092 19654
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18156 18970 18184 19790
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17958 18864 18014 18873
rect 17604 18822 17724 18850
rect 17696 18630 17724 18822
rect 17958 18799 18014 18808
rect 18052 18828 18104 18834
rect 17972 18766 18000 18799
rect 18052 18770 18104 18776
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17707 18524 18015 18533
rect 17707 18522 17713 18524
rect 17769 18522 17793 18524
rect 17849 18522 17873 18524
rect 17929 18522 17953 18524
rect 18009 18522 18015 18524
rect 17769 18470 17771 18522
rect 17951 18470 17953 18522
rect 17707 18468 17713 18470
rect 17769 18468 17793 18470
rect 17849 18468 17873 18470
rect 17929 18468 17953 18470
rect 18009 18468 18015 18470
rect 17707 18459 18015 18468
rect 17707 17436 18015 17445
rect 17707 17434 17713 17436
rect 17769 17434 17793 17436
rect 17849 17434 17873 17436
rect 17929 17434 17953 17436
rect 18009 17434 18015 17436
rect 17769 17382 17771 17434
rect 17951 17382 17953 17434
rect 17707 17380 17713 17382
rect 17769 17380 17793 17382
rect 17849 17380 17873 17382
rect 17929 17380 17953 17382
rect 18009 17380 18015 17382
rect 17707 17371 18015 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16794 18000 17206
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18064 16454 18092 18770
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17604 16182 17632 16390
rect 17707 16348 18015 16357
rect 17707 16346 17713 16348
rect 17769 16346 17793 16348
rect 17849 16346 17873 16348
rect 17929 16346 17953 16348
rect 18009 16346 18015 16348
rect 17769 16294 17771 16346
rect 17951 16294 17953 16346
rect 17707 16292 17713 16294
rect 17769 16292 17793 16294
rect 17849 16292 17873 16294
rect 17929 16292 17953 16294
rect 18009 16292 18015 16294
rect 17707 16283 18015 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17682 16144 17738 16153
rect 17682 16079 17738 16088
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17696 15416 17724 16079
rect 17972 15570 18000 16186
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18064 15638 18092 16050
rect 18156 16046 18184 17614
rect 18248 17202 18276 19910
rect 18800 19854 18828 20470
rect 19156 20392 19208 20398
rect 25516 20369 25544 26318
rect 26160 25945 26188 26386
rect 26146 25936 26202 25945
rect 26146 25871 26202 25880
rect 19156 20334 19208 20340
rect 25502 20360 25558 20369
rect 19168 19854 19196 20334
rect 25502 20295 25558 20304
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18340 18630 18368 19722
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18616 18766 18644 19110
rect 18800 18766 18828 19790
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18892 18970 18920 19382
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18086 18368 18566
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18800 17241 18828 18702
rect 18984 18426 19012 19790
rect 19168 19514 19196 19790
rect 19536 19514 19564 19858
rect 19996 19786 20024 20198
rect 23486 20156 23794 20165
rect 23486 20154 23492 20156
rect 23548 20154 23572 20156
rect 23628 20154 23652 20156
rect 23708 20154 23732 20156
rect 23788 20154 23794 20156
rect 23548 20102 23550 20154
rect 23730 20102 23732 20154
rect 23486 20100 23492 20102
rect 23548 20100 23572 20102
rect 23628 20100 23652 20102
rect 23708 20100 23732 20102
rect 23788 20100 23794 20102
rect 23486 20091 23794 20100
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18786 17232 18842 17241
rect 18236 17196 18288 17202
rect 18786 17167 18842 17176
rect 18236 17138 18288 17144
rect 19076 17134 19104 17478
rect 19168 17270 19196 19450
rect 19536 18766 19564 19450
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 20088 18970 20116 19246
rect 20456 18970 20484 19382
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 18358 19472 18566
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19352 17338 19380 18090
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16590 18276 16934
rect 18340 16590 18368 17002
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18432 16658 18460 16730
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18248 16114 18276 16526
rect 18340 16454 18368 16526
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 16182 18368 16390
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18418 16144 18474 16153
rect 18236 16108 18288 16114
rect 18418 16079 18420 16088
rect 18236 16050 18288 16056
rect 18472 16079 18474 16088
rect 18420 16050 18472 16056
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17604 15388 17724 15416
rect 18052 15428 18104 15434
rect 17604 15144 17632 15388
rect 18052 15370 18104 15376
rect 17707 15260 18015 15269
rect 17707 15258 17713 15260
rect 17769 15258 17793 15260
rect 17849 15258 17873 15260
rect 17929 15258 17953 15260
rect 18009 15258 18015 15260
rect 17769 15206 17771 15258
rect 17951 15206 17953 15258
rect 17707 15204 17713 15206
rect 17769 15204 17793 15206
rect 17849 15204 17873 15206
rect 17929 15204 17953 15206
rect 18009 15204 18015 15206
rect 17707 15195 18015 15204
rect 17604 15116 17724 15144
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 13870 17540 14214
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 17047 13628 17355 13637
rect 17047 13626 17053 13628
rect 17109 13626 17133 13628
rect 17189 13626 17213 13628
rect 17269 13626 17293 13628
rect 17349 13626 17355 13628
rect 17109 13574 17111 13626
rect 17291 13574 17293 13626
rect 17047 13572 17053 13574
rect 17109 13572 17133 13574
rect 17189 13572 17213 13574
rect 17269 13572 17293 13574
rect 17349 13572 17355 13574
rect 17047 13563 17355 13572
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12442 16988 13194
rect 17512 12986 17540 13398
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17047 12540 17355 12549
rect 17047 12538 17053 12540
rect 17109 12538 17133 12540
rect 17189 12538 17213 12540
rect 17269 12538 17293 12540
rect 17349 12538 17355 12540
rect 17109 12486 17111 12538
rect 17291 12486 17293 12538
rect 17047 12484 17053 12486
rect 17109 12484 17133 12486
rect 17189 12484 17213 12486
rect 17269 12484 17293 12486
rect 17349 12484 17355 12486
rect 17047 12475 17355 12484
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17604 12306 17632 14826
rect 17696 14618 17724 15116
rect 18064 14906 18092 15370
rect 18248 15162 18276 16050
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18340 15366 18368 15574
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17972 14878 18092 14906
rect 17972 14618 18000 14878
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 14521 18000 14554
rect 17958 14512 18014 14521
rect 18064 14482 18092 14758
rect 17958 14447 18014 14456
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17707 14172 18015 14181
rect 17707 14170 17713 14172
rect 17769 14170 17793 14172
rect 17849 14170 17873 14172
rect 17929 14170 17953 14172
rect 18009 14170 18015 14172
rect 17769 14118 17771 14170
rect 17951 14118 17953 14170
rect 17707 14116 17713 14118
rect 17769 14116 17793 14118
rect 17849 14116 17873 14118
rect 17929 14116 17953 14118
rect 18009 14116 18015 14118
rect 17707 14107 18015 14116
rect 18064 13802 18092 14418
rect 18156 14074 18184 14962
rect 18340 14822 18368 15302
rect 18432 14958 18460 15438
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18328 14816 18380 14822
rect 18380 14776 18460 14804
rect 18328 14758 18380 14764
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18340 14521 18368 14554
rect 18432 14550 18460 14776
rect 18420 14544 18472 14550
rect 18326 14512 18382 14521
rect 18420 14486 18472 14492
rect 18524 14482 18552 16526
rect 18326 14447 18382 14456
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18328 14386 18380 14392
rect 18708 14346 18736 16730
rect 18800 16658 18828 17002
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18984 16114 19012 16662
rect 19168 16130 19196 17206
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 16726 19288 16934
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19076 16114 19196 16130
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 19064 16108 19196 16114
rect 19116 16102 19196 16108
rect 19064 16050 19116 16056
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15706 19380 15982
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18800 15026 18828 15506
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 19076 14958 19104 15370
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 18892 14618 18920 14758
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18786 14376 18842 14385
rect 18328 14328 18380 14334
rect 18696 14340 18748 14346
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18156 13410 18184 14010
rect 18340 14006 18368 14328
rect 18786 14311 18842 14320
rect 18696 14282 18748 14288
rect 18708 14074 18736 14282
rect 18800 14278 18828 14311
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18064 13394 18184 13410
rect 18052 13388 18184 13394
rect 18104 13382 18184 13388
rect 18052 13330 18104 13336
rect 18340 13326 18368 13806
rect 18616 13394 18644 13874
rect 18892 13734 18920 14554
rect 19064 14544 19116 14550
rect 19062 14512 19064 14521
rect 19116 14512 19118 14521
rect 18972 14476 19024 14482
rect 19062 14447 19118 14456
rect 18972 14418 19024 14424
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18892 13530 18920 13670
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18144 13320 18196 13326
rect 18328 13320 18380 13326
rect 18196 13280 18276 13308
rect 18144 13262 18196 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 17707 13084 18015 13093
rect 17707 13082 17713 13084
rect 17769 13082 17793 13084
rect 17849 13082 17873 13084
rect 17929 13082 17953 13084
rect 18009 13082 18015 13084
rect 17769 13030 17771 13082
rect 17951 13030 17953 13082
rect 17707 13028 17713 13030
rect 17769 13028 17793 13030
rect 17849 13028 17873 13030
rect 17929 13028 17953 13030
rect 18009 13028 18015 13030
rect 17707 13019 18015 13028
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 18064 12238 18092 12786
rect 18156 12782 18184 13126
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16776 11898 16804 12106
rect 18248 12102 18276 13280
rect 18328 13262 18380 13268
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12918 18736 13262
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18984 12832 19012 14418
rect 19076 14414 19104 14447
rect 19168 14414 19196 14758
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19260 13394 19288 14894
rect 19444 14278 19472 16730
rect 19812 16454 19840 18770
rect 21008 18426 21036 19654
rect 24146 19612 24454 19621
rect 24146 19610 24152 19612
rect 24208 19610 24232 19612
rect 24288 19610 24312 19612
rect 24368 19610 24392 19612
rect 24448 19610 24454 19612
rect 24208 19558 24210 19610
rect 24390 19558 24392 19610
rect 24146 19556 24152 19558
rect 24208 19556 24232 19558
rect 24288 19556 24312 19558
rect 24368 19556 24392 19558
rect 24448 19556 24454 19558
rect 24146 19547 24454 19556
rect 23486 19068 23794 19077
rect 23486 19066 23492 19068
rect 23548 19066 23572 19068
rect 23628 19066 23652 19068
rect 23708 19066 23732 19068
rect 23788 19066 23794 19068
rect 23548 19014 23550 19066
rect 23730 19014 23732 19066
rect 23486 19012 23492 19014
rect 23548 19012 23572 19014
rect 23628 19012 23652 19014
rect 23708 19012 23732 19014
rect 23788 19012 23794 19014
rect 23486 19003 23794 19012
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26528 18601 26556 18702
rect 26514 18592 26570 18601
rect 24146 18524 24454 18533
rect 26514 18527 26570 18536
rect 24146 18522 24152 18524
rect 24208 18522 24232 18524
rect 24288 18522 24312 18524
rect 24368 18522 24392 18524
rect 24448 18522 24454 18524
rect 24208 18470 24210 18522
rect 24390 18470 24392 18522
rect 24146 18468 24152 18470
rect 24208 18468 24232 18470
rect 24288 18468 24312 18470
rect 24368 18468 24392 18470
rect 24448 18468 24454 18470
rect 24146 18459 24454 18468
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 23486 17980 23794 17989
rect 23486 17978 23492 17980
rect 23548 17978 23572 17980
rect 23628 17978 23652 17980
rect 23708 17978 23732 17980
rect 23788 17978 23794 17980
rect 23548 17926 23550 17978
rect 23730 17926 23732 17978
rect 23486 17924 23492 17926
rect 23548 17924 23572 17926
rect 23628 17924 23652 17926
rect 23708 17924 23732 17926
rect 23788 17924 23794 17926
rect 23486 17915 23794 17924
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 16182 20392 16390
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19536 14618 19564 14894
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19812 14482 19840 15302
rect 19904 15162 19932 15438
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19904 14550 19932 15098
rect 20732 14822 20760 15982
rect 20824 15502 20852 17138
rect 21652 16658 21680 17546
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 16182 21404 16526
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15570 21036 15846
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19812 13870 19840 14418
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 20640 13394 20668 14554
rect 20732 14482 20760 14758
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 19064 12844 19116 12850
rect 18984 12804 19064 12832
rect 19064 12786 19116 12792
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16854 11792 16910 11801
rect 17328 11762 17356 12038
rect 17707 11996 18015 12005
rect 17707 11994 17713 11996
rect 17769 11994 17793 11996
rect 17849 11994 17873 11996
rect 17929 11994 17953 11996
rect 18009 11994 18015 11996
rect 17769 11942 17771 11994
rect 17951 11942 17953 11994
rect 17707 11940 17713 11942
rect 17769 11940 17793 11942
rect 17849 11940 17873 11942
rect 17929 11940 17953 11942
rect 18009 11940 18015 11942
rect 17707 11931 18015 11940
rect 18064 11898 18092 12038
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 16854 11727 16856 11736
rect 16908 11727 16910 11736
rect 17316 11756 17368 11762
rect 16856 11698 16908 11704
rect 17316 11698 17368 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 17047 11452 17355 11461
rect 17047 11450 17053 11452
rect 17109 11450 17133 11452
rect 17189 11450 17213 11452
rect 17269 11450 17293 11452
rect 17349 11450 17355 11452
rect 17109 11398 17111 11450
rect 17291 11398 17293 11450
rect 17047 11396 17053 11398
rect 17109 11396 17133 11398
rect 17189 11396 17213 11398
rect 17269 11396 17293 11398
rect 17349 11396 17355 11398
rect 17047 11387 17355 11396
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 18432 11150 18460 12582
rect 18524 11150 18552 12582
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18800 11801 18828 12174
rect 19076 12170 19104 12242
rect 19260 12238 19288 13330
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 12986 20116 13194
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20640 12782 20668 13330
rect 20824 12850 20852 15438
rect 21376 15434 21404 16118
rect 21652 15706 21680 16458
rect 21836 16114 21864 17614
rect 24146 17436 24454 17445
rect 24146 17434 24152 17436
rect 24208 17434 24232 17436
rect 24288 17434 24312 17436
rect 24368 17434 24392 17436
rect 24448 17434 24454 17436
rect 24208 17382 24210 17434
rect 24390 17382 24392 17434
rect 24146 17380 24152 17382
rect 24208 17380 24232 17382
rect 24288 17380 24312 17382
rect 24368 17380 24392 17382
rect 24448 17380 24454 17382
rect 24146 17371 24454 17380
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21836 15706 21864 16050
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22112 15502 22140 16934
rect 22940 16794 22968 17138
rect 23032 16794 23060 17138
rect 23486 16892 23794 16901
rect 23486 16890 23492 16892
rect 23548 16890 23572 16892
rect 23628 16890 23652 16892
rect 23708 16890 23732 16892
rect 23788 16890 23794 16892
rect 23548 16838 23550 16890
rect 23730 16838 23732 16890
rect 23486 16836 23492 16838
rect 23548 16836 23572 16838
rect 23628 16836 23652 16838
rect 23708 16836 23732 16838
rect 23788 16836 23794 16838
rect 23486 16827 23794 16836
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22296 15638 22324 16458
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 16182 22508 16390
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22572 15910 22600 16526
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20916 15094 20944 15302
rect 21008 15162 21036 15370
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20994 13288 21050 13297
rect 20994 13223 21050 13232
rect 21008 12986 21036 13223
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11830 18920 12038
rect 18880 11824 18932 11830
rect 18786 11792 18842 11801
rect 18880 11766 18932 11772
rect 18786 11727 18842 11736
rect 19260 11218 19288 12174
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19444 11762 19472 12106
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17707 10908 18015 10917
rect 17707 10906 17713 10908
rect 17769 10906 17793 10908
rect 17849 10906 17873 10908
rect 17929 10906 17953 10908
rect 18009 10906 18015 10908
rect 17769 10854 17771 10906
rect 17951 10854 17953 10906
rect 17707 10852 17713 10854
rect 17769 10852 17793 10854
rect 17849 10852 17873 10854
rect 17929 10852 17953 10854
rect 18009 10852 18015 10854
rect 17707 10843 18015 10852
rect 19444 10674 19472 11698
rect 19536 11354 19564 12106
rect 19996 11762 20024 12718
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12306 20852 12650
rect 20916 12442 20944 12786
rect 21008 12714 21036 12922
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20088 11898 20116 12106
rect 20916 11898 20944 12378
rect 21376 12374 21404 15370
rect 22848 15366 22876 15982
rect 22940 15366 22968 16730
rect 23848 16720 23900 16726
rect 23848 16662 23900 16668
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23216 15910 23244 16390
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22848 15026 22876 15302
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 23216 14890 23244 15846
rect 23400 15502 23428 15846
rect 23486 15804 23794 15813
rect 23486 15802 23492 15804
rect 23548 15802 23572 15804
rect 23628 15802 23652 15804
rect 23708 15802 23732 15804
rect 23788 15802 23794 15804
rect 23548 15750 23550 15802
rect 23730 15750 23732 15802
rect 23486 15748 23492 15750
rect 23548 15748 23572 15750
rect 23628 15748 23652 15750
rect 23708 15748 23732 15750
rect 23788 15748 23794 15750
rect 23486 15739 23794 15748
rect 23388 15496 23440 15502
rect 23860 15484 23888 16662
rect 24032 16584 24084 16590
rect 23952 16532 24032 16538
rect 23952 16526 24084 16532
rect 23952 16510 24072 16526
rect 23952 16250 23980 16510
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 24044 16114 24072 16390
rect 24146 16348 24454 16357
rect 24146 16346 24152 16348
rect 24208 16346 24232 16348
rect 24288 16346 24312 16348
rect 24368 16346 24392 16348
rect 24448 16346 24454 16348
rect 24208 16294 24210 16346
rect 24390 16294 24392 16346
rect 24146 16292 24152 16294
rect 24208 16292 24232 16294
rect 24288 16292 24312 16294
rect 24368 16292 24392 16294
rect 24448 16292 24454 16294
rect 24146 16283 24454 16292
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24492 15972 24544 15978
rect 24492 15914 24544 15920
rect 24032 15496 24084 15502
rect 23860 15456 24032 15484
rect 23388 15438 23440 15444
rect 24032 15438 24084 15444
rect 24044 15094 24072 15438
rect 24146 15260 24454 15269
rect 24146 15258 24152 15260
rect 24208 15258 24232 15260
rect 24288 15258 24312 15260
rect 24368 15258 24392 15260
rect 24448 15258 24454 15260
rect 24208 15206 24210 15258
rect 24390 15206 24392 15258
rect 24146 15204 24152 15206
rect 24208 15204 24232 15206
rect 24288 15204 24312 15206
rect 24368 15204 24392 15206
rect 24448 15204 24454 15206
rect 24146 15195 24454 15204
rect 24504 15162 24532 15914
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 22480 14414 22508 14826
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 13938 22232 14214
rect 22572 14074 22600 14350
rect 22664 14074 22692 14350
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22756 13938 22784 14758
rect 23486 14716 23794 14725
rect 23486 14714 23492 14716
rect 23548 14714 23572 14716
rect 23628 14714 23652 14716
rect 23708 14714 23732 14716
rect 23788 14714 23794 14716
rect 23548 14662 23550 14714
rect 23730 14662 23732 14714
rect 23486 14660 23492 14662
rect 23548 14660 23572 14662
rect 23628 14660 23652 14662
rect 23708 14660 23732 14662
rect 23788 14660 23794 14662
rect 23486 14651 23794 14660
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 13530 22140 13806
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19628 10810 19656 11018
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 17047 10364 17355 10373
rect 17047 10362 17053 10364
rect 17109 10362 17133 10364
rect 17189 10362 17213 10364
rect 17269 10362 17293 10364
rect 17349 10362 17355 10364
rect 17109 10310 17111 10362
rect 17291 10310 17293 10362
rect 17047 10308 17053 10310
rect 17109 10308 17133 10310
rect 17189 10308 17213 10310
rect 17269 10308 17293 10310
rect 17349 10308 17355 10310
rect 17047 10299 17355 10308
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 17707 9820 18015 9829
rect 17707 9818 17713 9820
rect 17769 9818 17793 9820
rect 17849 9818 17873 9820
rect 17929 9818 17953 9820
rect 18009 9818 18015 9820
rect 17769 9766 17771 9818
rect 17951 9766 17953 9818
rect 17707 9764 17713 9766
rect 17769 9764 17793 9766
rect 17849 9764 17873 9766
rect 17929 9764 17953 9766
rect 18009 9764 18015 9766
rect 17707 9755 18015 9764
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16684 9178 16712 9590
rect 19444 9586 19472 9998
rect 21376 9994 21404 12310
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21468 11626 21496 12106
rect 21652 11830 21680 12378
rect 21836 12238 21864 12582
rect 22020 12442 22048 12786
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21744 11558 21772 11766
rect 22008 11756 22060 11762
rect 22112 11744 22140 13466
rect 22388 11830 22416 13874
rect 22848 13530 22876 14350
rect 22940 13870 22968 14350
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22940 13326 22968 13806
rect 23032 13802 23060 13874
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23216 13462 23244 14350
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23768 13938 23796 14214
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23308 13394 23336 13874
rect 23492 13818 23520 13874
rect 23400 13790 23520 13818
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22848 12442 22876 13262
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 23032 12306 23060 13330
rect 23400 13326 23428 13790
rect 23486 13628 23794 13637
rect 23486 13626 23492 13628
rect 23548 13626 23572 13628
rect 23628 13626 23652 13628
rect 23708 13626 23732 13628
rect 23788 13626 23794 13628
rect 23548 13574 23550 13626
rect 23730 13574 23732 13626
rect 23486 13572 23492 13574
rect 23548 13572 23572 13574
rect 23628 13572 23652 13574
rect 23708 13572 23732 13574
rect 23788 13572 23794 13574
rect 23486 13563 23794 13572
rect 23860 13462 23888 14214
rect 23952 13462 23980 14418
rect 24044 14056 24072 15030
rect 24504 14958 24532 15098
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 24136 14346 24164 14826
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 14414 24256 14758
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24124 14340 24176 14346
rect 24124 14282 24176 14288
rect 24146 14172 24454 14181
rect 24146 14170 24152 14172
rect 24208 14170 24232 14172
rect 24288 14170 24312 14172
rect 24368 14170 24392 14172
rect 24448 14170 24454 14172
rect 24208 14118 24210 14170
rect 24390 14118 24392 14170
rect 24146 14116 24152 14118
rect 24208 14116 24232 14118
rect 24288 14116 24312 14118
rect 24368 14116 24392 14118
rect 24448 14116 24454 14118
rect 24146 14107 24454 14116
rect 24044 14028 24164 14056
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 24044 13326 24072 13670
rect 24136 13530 24164 14028
rect 24504 14006 24532 14894
rect 24596 14890 24624 16050
rect 25056 15162 25084 16050
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 25148 15502 25176 15846
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25884 14958 25912 15302
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24596 14498 24624 14826
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24596 14470 24808 14498
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24596 13394 24624 14350
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24780 13818 24808 14470
rect 24872 14074 24900 14554
rect 25056 14346 25084 14894
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24584 13388 24636 13394
rect 24504 13348 24584 13376
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23952 12986 23980 13262
rect 24146 13084 24454 13093
rect 24146 13082 24152 13084
rect 24208 13082 24232 13084
rect 24288 13082 24312 13084
rect 24368 13082 24392 13084
rect 24448 13082 24454 13084
rect 24208 13030 24210 13082
rect 24390 13030 24392 13082
rect 24146 13028 24152 13030
rect 24208 13028 24232 13030
rect 24288 13028 24312 13030
rect 24368 13028 24392 13030
rect 24448 13028 24454 13030
rect 24146 13019 24454 13028
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23486 12540 23794 12549
rect 23486 12538 23492 12540
rect 23548 12538 23572 12540
rect 23628 12538 23652 12540
rect 23708 12538 23732 12540
rect 23788 12538 23794 12540
rect 23548 12486 23550 12538
rect 23730 12486 23732 12538
rect 23486 12484 23492 12486
rect 23548 12484 23572 12486
rect 23628 12484 23652 12486
rect 23708 12484 23732 12486
rect 23788 12484 23794 12486
rect 23486 12475 23794 12484
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22664 11762 22692 12038
rect 23032 11762 23060 12242
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 22192 11756 22244 11762
rect 22112 11716 22192 11744
rect 22008 11698 22060 11704
rect 22192 11698 22244 11704
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21836 10742 21864 11562
rect 22020 11354 22048 11698
rect 22204 11354 22232 11698
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22204 11218 22232 11290
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22480 11150 22508 11698
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22940 11354 22968 11630
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22756 11150 22784 11290
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 21836 10266 21864 10678
rect 22112 10674 22140 11086
rect 22480 10826 22508 11086
rect 23032 11082 23060 11698
rect 23124 11098 23152 12174
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23216 11354 23244 11698
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23400 11286 23428 12310
rect 24146 11996 24454 12005
rect 24146 11994 24152 11996
rect 24208 11994 24232 11996
rect 24288 11994 24312 11996
rect 24368 11994 24392 11996
rect 24448 11994 24454 11996
rect 24208 11942 24210 11994
rect 24390 11942 24392 11994
rect 24146 11940 24152 11942
rect 24208 11940 24232 11942
rect 24288 11940 24312 11942
rect 24368 11940 24392 11942
rect 24448 11940 24454 11942
rect 24146 11931 24454 11940
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23486 11452 23794 11461
rect 23486 11450 23492 11452
rect 23548 11450 23572 11452
rect 23628 11450 23652 11452
rect 23708 11450 23732 11452
rect 23788 11450 23794 11452
rect 23548 11398 23550 11450
rect 23730 11398 23732 11450
rect 23486 11396 23492 11398
rect 23548 11396 23572 11398
rect 23628 11396 23652 11398
rect 23708 11396 23732 11398
rect 23788 11396 23794 11398
rect 23486 11387 23794 11396
rect 23952 11354 23980 11494
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23124 11082 23244 11098
rect 23020 11076 23072 11082
rect 23124 11076 23256 11082
rect 23124 11070 23204 11076
rect 23020 11018 23072 11024
rect 23204 11018 23256 11024
rect 22480 10810 22600 10826
rect 22480 10804 22612 10810
rect 22480 10798 22560 10804
rect 22560 10746 22612 10752
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22204 10266 22232 10406
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22296 10248 22324 10406
rect 22376 10260 22428 10266
rect 22296 10220 22376 10248
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21364 9988 21416 9994
rect 21364 9930 21416 9936
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21284 9722 21312 9930
rect 21928 9722 21956 9930
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9722 22140 9862
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22296 9602 22324 10220
rect 22376 10202 22428 10208
rect 22756 10130 22784 10406
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22940 9654 22968 10610
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 22112 9574 22324 9602
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 23032 9586 23060 9862
rect 23216 9654 23244 11018
rect 24146 10908 24454 10917
rect 24146 10906 24152 10908
rect 24208 10906 24232 10908
rect 24288 10906 24312 10908
rect 24368 10906 24392 10908
rect 24448 10906 24454 10908
rect 24208 10854 24210 10906
rect 24390 10854 24392 10906
rect 24146 10852 24152 10854
rect 24208 10852 24232 10854
rect 24288 10852 24312 10854
rect 24368 10852 24392 10854
rect 24448 10852 24454 10854
rect 24146 10843 24454 10852
rect 24504 10674 24532 13348
rect 24584 13330 24636 13336
rect 24688 12986 24716 13806
rect 24780 13790 24900 13818
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24872 12850 24900 13790
rect 25056 13734 25084 14282
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24964 12986 24992 13194
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25332 12850 25360 14010
rect 25976 13938 26004 14214
rect 26436 14074 26464 14962
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 23486 10364 23794 10373
rect 23486 10362 23492 10364
rect 23548 10362 23572 10364
rect 23628 10362 23652 10364
rect 23708 10362 23732 10364
rect 23788 10362 23794 10364
rect 23548 10310 23550 10362
rect 23730 10310 23732 10362
rect 23486 10308 23492 10310
rect 23548 10308 23572 10310
rect 23628 10308 23652 10310
rect 23708 10308 23732 10310
rect 23788 10308 23794 10310
rect 23486 10299 23794 10308
rect 24044 9722 24072 10406
rect 24504 10130 24532 10610
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24146 9820 24454 9829
rect 24146 9818 24152 9820
rect 24208 9818 24232 9820
rect 24288 9818 24312 9820
rect 24368 9818 24392 9820
rect 24448 9818 24454 9820
rect 24208 9766 24210 9818
rect 24390 9766 24392 9818
rect 24146 9764 24152 9766
rect 24208 9764 24232 9766
rect 24288 9764 24312 9766
rect 24368 9764 24392 9766
rect 24448 9764 24454 9766
rect 24146 9755 24454 9764
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23020 9580 23072 9586
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16776 8974 16804 9318
rect 17047 9276 17355 9285
rect 17047 9274 17053 9276
rect 17109 9274 17133 9276
rect 17189 9274 17213 9276
rect 17269 9274 17293 9276
rect 17349 9274 17355 9276
rect 17109 9222 17111 9274
rect 17291 9222 17293 9274
rect 17047 9220 17053 9222
rect 17109 9220 17133 9222
rect 17189 9220 17213 9222
rect 17269 9220 17293 9222
rect 17349 9220 17355 9222
rect 17047 9211 17355 9220
rect 18156 9178 18184 9454
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18064 9042 18276 9058
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 18052 9036 18288 9042
rect 18104 9030 18236 9036
rect 18052 8978 18104 8984
rect 18236 8978 18288 8984
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 17144 8498 17172 8978
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 8378 17172 8434
rect 16960 8350 17172 8378
rect 17236 8362 17264 8910
rect 18432 8906 18460 9114
rect 19444 9110 19472 9522
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 17707 8732 18015 8741
rect 17707 8730 17713 8732
rect 17769 8730 17793 8732
rect 17849 8730 17873 8732
rect 17929 8730 17953 8732
rect 18009 8730 18015 8732
rect 17769 8678 17771 8730
rect 17951 8678 17953 8730
rect 17707 8676 17713 8678
rect 17769 8676 17793 8678
rect 17849 8676 17873 8678
rect 17929 8676 17953 8678
rect 18009 8676 18015 8678
rect 17707 8667 18015 8676
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17328 8430 17356 8570
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17224 8356 17276 8362
rect 16960 7546 16988 8350
rect 17224 8298 17276 8304
rect 17047 8188 17355 8197
rect 17047 8186 17053 8188
rect 17109 8186 17133 8188
rect 17189 8186 17213 8188
rect 17269 8186 17293 8188
rect 17349 8186 17355 8188
rect 17109 8134 17111 8186
rect 17291 8134 17293 8186
rect 17047 8132 17053 8134
rect 17109 8132 17133 8134
rect 17189 8132 17213 8134
rect 17269 8132 17293 8134
rect 17349 8132 17355 8134
rect 17047 8123 17355 8132
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16960 7274 16988 7346
rect 17052 7313 17080 7346
rect 17038 7304 17094 7313
rect 16948 7268 17000 7274
rect 17038 7239 17094 7248
rect 16948 7210 17000 7216
rect 17047 7100 17355 7109
rect 17047 7098 17053 7100
rect 17109 7098 17133 7100
rect 17189 7098 17213 7100
rect 17269 7098 17293 7100
rect 17349 7098 17355 7100
rect 17109 7046 17111 7098
rect 17291 7046 17293 7098
rect 17047 7044 17053 7046
rect 17109 7044 17133 7046
rect 17189 7044 17213 7046
rect 17269 7044 17293 7046
rect 17349 7044 17355 7046
rect 17047 7035 17355 7044
rect 17420 6866 17448 8366
rect 17972 8362 18000 8434
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17707 7644 18015 7653
rect 17707 7642 17713 7644
rect 17769 7642 17793 7644
rect 17849 7642 17873 7644
rect 17929 7642 17953 7644
rect 18009 7642 18015 7644
rect 17769 7590 17771 7642
rect 17951 7590 17953 7642
rect 17707 7588 17713 7590
rect 17769 7588 17793 7590
rect 17849 7588 17873 7590
rect 17929 7588 17953 7590
rect 18009 7588 18015 7590
rect 17707 7579 18015 7588
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 16684 5710 16712 6802
rect 17696 6798 17724 7346
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 16960 6458 16988 6666
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17420 6390 17448 6666
rect 18064 6662 18092 8298
rect 18156 8090 18184 8774
rect 18340 8634 18368 8774
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18340 8090 18368 8434
rect 18432 8294 18460 8842
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8566 18552 8774
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18708 8498 18736 8842
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18708 7886 18736 8298
rect 18984 7886 19012 8366
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7410 18184 7686
rect 18800 7546 18828 7822
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17707 6556 18015 6565
rect 17707 6554 17713 6556
rect 17769 6554 17793 6556
rect 17849 6554 17873 6556
rect 17929 6554 17953 6556
rect 18009 6554 18015 6556
rect 17769 6502 17771 6554
rect 17951 6502 17953 6554
rect 17707 6500 17713 6502
rect 17769 6500 17793 6502
rect 17849 6500 17873 6502
rect 17929 6500 17953 6502
rect 18009 6500 18015 6502
rect 17707 6491 18015 6500
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17047 6012 17355 6021
rect 17047 6010 17053 6012
rect 17109 6010 17133 6012
rect 17189 6010 17213 6012
rect 17269 6010 17293 6012
rect 17349 6010 17355 6012
rect 17109 5958 17111 6010
rect 17291 5958 17293 6010
rect 17047 5956 17053 5958
rect 17109 5956 17133 5958
rect 17189 5956 17213 5958
rect 17269 5956 17293 5958
rect 17349 5956 17355 5958
rect 17047 5947 17355 5956
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 18248 5574 18276 7346
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18892 6798 18920 7142
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18708 6322 18736 6734
rect 18892 6390 18920 6734
rect 19076 6662 19104 8366
rect 19260 7886 19288 9046
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8022 19380 8774
rect 19444 8498 19472 9046
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19260 7410 19288 7822
rect 19444 7546 19472 8434
rect 19536 7886 19564 8570
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19812 8090 19840 8366
rect 19984 8288 20036 8294
rect 19904 8248 19984 8276
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19904 7954 19932 8248
rect 19984 8230 20036 8236
rect 20364 8090 20392 8842
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 8566 20576 8774
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 19996 7954 20116 7970
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19996 7948 20128 7954
rect 19996 7942 20076 7948
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19536 7342 19564 7822
rect 19800 7812 19852 7818
rect 19800 7754 19852 7760
rect 19812 7546 19840 7754
rect 19904 7750 19932 7890
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19996 7478 20024 7942
rect 20076 7890 20128 7896
rect 20260 7880 20312 7886
rect 20180 7840 20260 7868
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 17707 5468 18015 5477
rect 17707 5466 17713 5468
rect 17769 5466 17793 5468
rect 17849 5466 17873 5468
rect 17929 5466 17953 5468
rect 18009 5466 18015 5468
rect 17769 5414 17771 5466
rect 17951 5414 17953 5466
rect 17707 5412 17713 5414
rect 17769 5412 17793 5414
rect 17849 5412 17873 5414
rect 17929 5412 17953 5414
rect 18009 5412 18015 5414
rect 17707 5403 18015 5412
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16592 4690 16620 5170
rect 18340 5166 18368 6190
rect 19168 5642 19196 6666
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 17047 4924 17355 4933
rect 17047 4922 17053 4924
rect 17109 4922 17133 4924
rect 17189 4922 17213 4924
rect 17269 4922 17293 4924
rect 17349 4922 17355 4924
rect 17109 4870 17111 4922
rect 17291 4870 17293 4922
rect 17047 4868 17053 4870
rect 17109 4868 17133 4870
rect 17189 4868 17213 4870
rect 17269 4868 17293 4870
rect 17349 4868 17355 4870
rect 17047 4859 17355 4868
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16592 4010 16620 4626
rect 16764 4616 16816 4622
rect 17052 4570 17080 4626
rect 16816 4564 17080 4570
rect 16764 4558 17080 4564
rect 16776 4542 17080 4558
rect 16948 4480 17000 4486
rect 16762 4448 16818 4457
rect 16948 4422 17000 4428
rect 16762 4383 16818 4392
rect 16776 4214 16804 4383
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3126 16896 3538
rect 16960 3126 16988 4422
rect 17052 4146 17080 4542
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17236 4146 17264 4422
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17420 4078 17448 4762
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 17707 4380 18015 4389
rect 17707 4378 17713 4380
rect 17769 4378 17793 4380
rect 17849 4378 17873 4380
rect 17929 4378 17953 4380
rect 18009 4378 18015 4380
rect 17769 4326 17771 4378
rect 17951 4326 17953 4378
rect 17707 4324 17713 4326
rect 17769 4324 17793 4326
rect 17849 4324 17873 4326
rect 17929 4324 17953 4326
rect 18009 4324 18015 4326
rect 17707 4315 18015 4324
rect 18064 4282 18092 4626
rect 18248 4554 18276 4694
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18156 4146 18184 4422
rect 18248 4146 18276 4490
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17408 4072 17460 4078
rect 17788 4049 17816 4082
rect 17408 4014 17460 4020
rect 17774 4040 17830 4049
rect 17328 3942 17356 4014
rect 17774 3975 17830 3984
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17047 3836 17355 3845
rect 17047 3834 17053 3836
rect 17109 3834 17133 3836
rect 17189 3834 17213 3836
rect 17269 3834 17293 3836
rect 17349 3834 17355 3836
rect 17109 3782 17111 3834
rect 17291 3782 17293 3834
rect 17047 3780 17053 3782
rect 17109 3780 17133 3782
rect 17189 3780 17213 3782
rect 17269 3780 17293 3782
rect 17349 3780 17355 3782
rect 17047 3771 17355 3780
rect 17696 3534 17724 3878
rect 18340 3534 18368 5102
rect 19168 4690 19196 5578
rect 19352 5370 19380 5782
rect 19536 5710 19564 7278
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19996 6662 20024 6734
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6322 20024 6598
rect 20088 6458 20116 7346
rect 20180 7274 20208 7840
rect 20260 7822 20312 7828
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20180 6934 20208 7210
rect 20168 6928 20220 6934
rect 20168 6870 20220 6876
rect 20180 6798 20208 6870
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5710 19656 6054
rect 20088 5846 20116 6394
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 20364 5778 20392 8026
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20456 7206 20484 7890
rect 20640 7834 20668 7890
rect 20548 7806 20668 7834
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5250 19472 5578
rect 19536 5574 19564 5646
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19352 5234 19472 5250
rect 19628 5234 19656 5646
rect 19340 5228 19472 5234
rect 19392 5222 19472 5228
rect 19340 5170 19392 5176
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18432 4146 18460 4558
rect 19168 4162 19196 4626
rect 19076 4146 19196 4162
rect 19260 4146 19288 4966
rect 19444 4690 19472 5222
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19996 4554 20024 4966
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 20456 4282 20484 7142
rect 20548 7002 20576 7806
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20640 7410 20668 7686
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20732 6186 20760 8434
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20824 7410 20852 7958
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7478 20944 7686
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 21008 7410 21036 7822
rect 21284 7546 21312 8842
rect 21744 8838 21772 9522
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21744 8498 21772 8774
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21652 7478 21680 8230
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20824 4826 20852 6258
rect 20916 6186 20944 7278
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 6866 21036 7142
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21100 6798 21128 7414
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 7002 21496 7142
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21468 6866 21496 6938
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21100 6390 21128 6734
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21468 6322 21496 6802
rect 21836 6322 21864 8978
rect 22112 8906 22140 9574
rect 23020 9522 23072 9528
rect 22744 9512 22796 9518
rect 23216 9466 23244 9590
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 22796 9460 23244 9466
rect 22744 9454 23244 9460
rect 22756 9438 23244 9454
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22204 9178 22232 9318
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22480 8634 22508 8842
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22664 8498 22692 8774
rect 22756 8634 22784 9438
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23216 9178 23244 9318
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23308 9110 23336 9522
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 9104 23348 9110
rect 23296 9046 23348 9052
rect 23400 8838 23428 9454
rect 23940 9444 23992 9450
rect 23940 9386 23992 9392
rect 23486 9276 23794 9285
rect 23486 9274 23492 9276
rect 23548 9274 23572 9276
rect 23628 9274 23652 9276
rect 23708 9274 23732 9276
rect 23788 9274 23794 9276
rect 23548 9222 23550 9274
rect 23730 9222 23732 9274
rect 23486 9220 23492 9222
rect 23548 9220 23572 9222
rect 23628 9220 23652 9222
rect 23708 9220 23732 9222
rect 23788 9220 23794 9222
rect 23486 9211 23794 9220
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 23676 8566 23704 8774
rect 23952 8634 23980 9386
rect 24044 9110 24072 9658
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24504 9042 24532 10066
rect 24596 10062 24624 11086
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 10810 24900 10950
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 25056 10470 25084 12786
rect 26252 12782 26280 13126
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 25792 11150 25820 11698
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25792 10810 25820 11086
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 9518 24624 9998
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24780 9586 24808 9930
rect 25056 9654 25084 10406
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9382 24624 9454
rect 25148 9382 25176 9862
rect 25332 9722 25360 9998
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 26068 9586 26096 9862
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24146 8732 24454 8741
rect 24146 8730 24152 8732
rect 24208 8730 24232 8732
rect 24288 8730 24312 8732
rect 24368 8730 24392 8732
rect 24448 8730 24454 8732
rect 24208 8678 24210 8730
rect 24390 8678 24392 8730
rect 24146 8676 24152 8678
rect 24208 8676 24232 8678
rect 24288 8676 24312 8678
rect 24368 8676 24392 8678
rect 24448 8676 24454 8678
rect 24146 8667 24454 8676
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 24504 8498 24532 8978
rect 26344 8974 26372 11494
rect 26528 11257 26556 11698
rect 26514 11248 26570 11257
rect 26514 11183 26570 11192
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 23486 8188 23794 8197
rect 23486 8186 23492 8188
rect 23548 8186 23572 8188
rect 23628 8186 23652 8188
rect 23708 8186 23732 8188
rect 23788 8186 23794 8188
rect 23548 8134 23550 8186
rect 23730 8134 23732 8186
rect 23486 8132 23492 8134
rect 23548 8132 23572 8134
rect 23628 8132 23652 8134
rect 23708 8132 23732 8134
rect 23788 8132 23794 8134
rect 23486 8123 23794 8132
rect 24146 7644 24454 7653
rect 24146 7642 24152 7644
rect 24208 7642 24232 7644
rect 24288 7642 24312 7644
rect 24368 7642 24392 7644
rect 24448 7642 24454 7644
rect 24208 7590 24210 7642
rect 24390 7590 24392 7642
rect 24146 7588 24152 7590
rect 24208 7588 24232 7590
rect 24288 7588 24312 7590
rect 24368 7588 24392 7590
rect 24448 7588 24454 7590
rect 24146 7579 24454 7588
rect 25700 7449 25728 8774
rect 25686 7440 25742 7449
rect 25686 7375 25742 7384
rect 23486 7100 23794 7109
rect 23486 7098 23492 7100
rect 23548 7098 23572 7100
rect 23628 7098 23652 7100
rect 23708 7098 23732 7100
rect 23788 7098 23794 7100
rect 23548 7046 23550 7098
rect 23730 7046 23732 7098
rect 23486 7044 23492 7046
rect 23548 7044 23572 7046
rect 23628 7044 23652 7046
rect 23708 7044 23732 7046
rect 23788 7044 23794 7046
rect 23486 7035 23794 7044
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21928 6458 21956 6666
rect 24146 6556 24454 6565
rect 24146 6554 24152 6556
rect 24208 6554 24232 6556
rect 24288 6554 24312 6556
rect 24368 6554 24392 6556
rect 24448 6554 24454 6556
rect 24208 6502 24210 6554
rect 24390 6502 24392 6554
rect 24146 6500 24152 6502
rect 24208 6500 24232 6502
rect 24288 6500 24312 6502
rect 24368 6500 24392 6502
rect 24448 6500 24454 6502
rect 24146 6491 24454 6500
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 21836 5166 21864 6258
rect 23486 6012 23794 6021
rect 23486 6010 23492 6012
rect 23548 6010 23572 6012
rect 23628 6010 23652 6012
rect 23708 6010 23732 6012
rect 23788 6010 23794 6012
rect 23548 5958 23550 6010
rect 23730 5958 23732 6010
rect 23486 5956 23492 5958
rect 23548 5956 23572 5958
rect 23628 5956 23652 5958
rect 23708 5956 23732 5958
rect 23788 5956 23794 5958
rect 23486 5947 23794 5956
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 24146 5468 24454 5477
rect 24146 5466 24152 5468
rect 24208 5466 24232 5468
rect 24288 5466 24312 5468
rect 24368 5466 24392 5468
rect 24448 5466 24454 5468
rect 24208 5414 24210 5466
rect 24390 5414 24392 5466
rect 24146 5412 24152 5414
rect 24208 5412 24232 5414
rect 24288 5412 24312 5414
rect 24368 5412 24392 5414
rect 24448 5412 24454 5414
rect 24146 5403 24454 5412
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20916 4146 20944 5102
rect 23486 4924 23794 4933
rect 23486 4922 23492 4924
rect 23548 4922 23572 4924
rect 23628 4922 23652 4924
rect 23708 4922 23732 4924
rect 23788 4922 23794 4924
rect 23548 4870 23550 4922
rect 23730 4870 23732 4922
rect 23486 4868 23492 4870
rect 23548 4868 23572 4870
rect 23628 4868 23652 4870
rect 23708 4868 23732 4870
rect 23788 4868 23794 4870
rect 23486 4859 23794 4868
rect 24146 4380 24454 4389
rect 24146 4378 24152 4380
rect 24208 4378 24232 4380
rect 24288 4378 24312 4380
rect 24368 4378 24392 4380
rect 24448 4378 24454 4380
rect 24208 4326 24210 4378
rect 24390 4326 24392 4378
rect 24146 4324 24152 4326
rect 24208 4324 24232 4326
rect 24288 4324 24312 4326
rect 24368 4324 24392 4326
rect 24448 4324 24454 4326
rect 24146 4315 24454 4324
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 19064 4140 19196 4146
rect 19116 4134 19196 4140
rect 19248 4140 19300 4146
rect 19064 4082 19116 4088
rect 19248 4082 19300 4088
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 17707 3292 18015 3301
rect 17707 3290 17713 3292
rect 17769 3290 17793 3292
rect 17849 3290 17873 3292
rect 17929 3290 17953 3292
rect 18009 3290 18015 3292
rect 17769 3238 17771 3290
rect 17951 3238 17953 3290
rect 17707 3236 17713 3238
rect 17769 3236 17793 3238
rect 17849 3236 17873 3238
rect 17929 3236 17953 3238
rect 18009 3236 18015 3238
rect 17707 3227 18015 3236
rect 18432 3194 18460 3946
rect 19076 3602 19104 4082
rect 26344 4010 26372 5646
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26332 4004 26384 4010
rect 26332 3946 26384 3952
rect 26528 3913 26556 4082
rect 26514 3904 26570 3913
rect 23486 3836 23794 3845
rect 26514 3839 26570 3848
rect 23486 3834 23492 3836
rect 23548 3834 23572 3836
rect 23628 3834 23652 3836
rect 23708 3834 23732 3836
rect 23788 3834 23794 3836
rect 23548 3782 23550 3834
rect 23730 3782 23732 3834
rect 23486 3780 23492 3782
rect 23548 3780 23572 3782
rect 23628 3780 23652 3782
rect 23708 3780 23732 3782
rect 23788 3780 23794 3782
rect 23486 3771 23794 3780
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18524 3126 18552 3334
rect 24146 3292 24454 3301
rect 24146 3290 24152 3292
rect 24208 3290 24232 3292
rect 24288 3290 24312 3292
rect 24368 3290 24392 3292
rect 24448 3290 24454 3292
rect 24208 3238 24210 3290
rect 24390 3238 24392 3290
rect 24146 3236 24152 3238
rect 24208 3236 24232 3238
rect 24288 3236 24312 3238
rect 24368 3236 24392 3238
rect 24448 3236 24454 3238
rect 24146 3227 24454 3236
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 17047 2748 17355 2757
rect 17047 2746 17053 2748
rect 17109 2746 17133 2748
rect 17189 2746 17213 2748
rect 17269 2746 17293 2748
rect 17349 2746 17355 2748
rect 17109 2694 17111 2746
rect 17291 2694 17293 2746
rect 17047 2692 17053 2694
rect 17109 2692 17133 2694
rect 17189 2692 17213 2694
rect 17269 2692 17293 2694
rect 17349 2692 17355 2694
rect 17047 2683 17355 2692
rect 23486 2748 23794 2757
rect 23486 2746 23492 2748
rect 23548 2746 23572 2748
rect 23628 2746 23652 2748
rect 23708 2746 23732 2748
rect 23788 2746 23794 2748
rect 23548 2694 23550 2746
rect 23730 2694 23732 2746
rect 23486 2692 23492 2694
rect 23548 2692 23572 2694
rect 23628 2692 23652 2694
rect 23708 2692 23732 2694
rect 23788 2692 23794 2694
rect 23486 2683 23794 2692
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 4829 2204 5137 2213
rect 4829 2202 4835 2204
rect 4891 2202 4915 2204
rect 4971 2202 4995 2204
rect 5051 2202 5075 2204
rect 5131 2202 5137 2204
rect 4891 2150 4893 2202
rect 5073 2150 5075 2202
rect 4829 2148 4835 2150
rect 4891 2148 4915 2150
rect 4971 2148 4995 2150
rect 5051 2148 5075 2150
rect 5131 2148 5137 2150
rect 4829 2139 5137 2148
rect 6012 800 6040 2314
rect 9968 800 9996 2314
rect 11268 2204 11576 2213
rect 11268 2202 11274 2204
rect 11330 2202 11354 2204
rect 11410 2202 11434 2204
rect 11490 2202 11514 2204
rect 11570 2202 11576 2204
rect 11330 2150 11332 2202
rect 11512 2150 11514 2202
rect 11268 2148 11274 2150
rect 11330 2148 11354 2150
rect 11410 2148 11434 2150
rect 11490 2148 11514 2150
rect 11570 2148 11576 2150
rect 11268 2139 11576 2148
rect 13924 800 13952 2314
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 17707 2204 18015 2213
rect 17707 2202 17713 2204
rect 17769 2202 17793 2204
rect 17849 2202 17873 2204
rect 17929 2202 17953 2204
rect 18009 2202 18015 2204
rect 17769 2150 17771 2202
rect 17951 2150 17953 2202
rect 17707 2148 17713 2150
rect 17769 2148 17793 2150
rect 17849 2148 17873 2150
rect 17929 2148 17953 2150
rect 18009 2148 18015 2150
rect 17707 2139 18015 2148
rect 18156 1442 18184 2246
rect 17880 1414 18184 1442
rect 17880 800 17908 1414
rect 21836 800 21864 2246
rect 24146 2204 24454 2213
rect 24146 2202 24152 2204
rect 24208 2202 24232 2204
rect 24288 2202 24312 2204
rect 24368 2202 24392 2204
rect 24448 2202 24454 2204
rect 24208 2150 24210 2202
rect 24390 2150 24392 2202
rect 24146 2148 24152 2150
rect 24208 2148 24232 2150
rect 24288 2148 24312 2150
rect 24368 2148 24392 2150
rect 24448 2148 24454 2150
rect 24146 2139 24454 2148
rect 25792 800 25820 2246
rect 2042 0 2098 800
rect 5998 0 6054 800
rect 9954 0 10010 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21822 0 21878 800
rect 25778 0 25834 800
<< via2 >>
rect 2226 28056 2282 28112
rect 938 23724 994 23760
rect 938 23704 940 23724
rect 940 23704 992 23724
rect 992 23704 994 23724
rect 938 21528 994 21584
rect 4175 27770 4231 27772
rect 4255 27770 4311 27772
rect 4335 27770 4391 27772
rect 4415 27770 4471 27772
rect 4175 27718 4221 27770
rect 4221 27718 4231 27770
rect 4255 27718 4285 27770
rect 4285 27718 4297 27770
rect 4297 27718 4311 27770
rect 4335 27718 4349 27770
rect 4349 27718 4361 27770
rect 4361 27718 4391 27770
rect 4415 27718 4425 27770
rect 4425 27718 4471 27770
rect 4175 27716 4231 27718
rect 4255 27716 4311 27718
rect 4335 27716 4391 27718
rect 4415 27716 4471 27718
rect 10614 27770 10670 27772
rect 10694 27770 10750 27772
rect 10774 27770 10830 27772
rect 10854 27770 10910 27772
rect 10614 27718 10660 27770
rect 10660 27718 10670 27770
rect 10694 27718 10724 27770
rect 10724 27718 10736 27770
rect 10736 27718 10750 27770
rect 10774 27718 10788 27770
rect 10788 27718 10800 27770
rect 10800 27718 10830 27770
rect 10854 27718 10864 27770
rect 10864 27718 10910 27770
rect 10614 27716 10670 27718
rect 10694 27716 10750 27718
rect 10774 27716 10830 27718
rect 10854 27716 10910 27718
rect 17053 27770 17109 27772
rect 17133 27770 17189 27772
rect 17213 27770 17269 27772
rect 17293 27770 17349 27772
rect 17053 27718 17099 27770
rect 17099 27718 17109 27770
rect 17133 27718 17163 27770
rect 17163 27718 17175 27770
rect 17175 27718 17189 27770
rect 17213 27718 17227 27770
rect 17227 27718 17239 27770
rect 17239 27718 17269 27770
rect 17293 27718 17303 27770
rect 17303 27718 17349 27770
rect 17053 27716 17109 27718
rect 17133 27716 17189 27718
rect 17213 27716 17269 27718
rect 17293 27716 17349 27718
rect 23492 27770 23548 27772
rect 23572 27770 23628 27772
rect 23652 27770 23708 27772
rect 23732 27770 23788 27772
rect 23492 27718 23538 27770
rect 23538 27718 23548 27770
rect 23572 27718 23602 27770
rect 23602 27718 23614 27770
rect 23614 27718 23628 27770
rect 23652 27718 23666 27770
rect 23666 27718 23678 27770
rect 23678 27718 23708 27770
rect 23732 27718 23742 27770
rect 23742 27718 23788 27770
rect 23492 27716 23548 27718
rect 23572 27716 23628 27718
rect 23652 27716 23708 27718
rect 23732 27716 23788 27718
rect 4835 27226 4891 27228
rect 4915 27226 4971 27228
rect 4995 27226 5051 27228
rect 5075 27226 5131 27228
rect 4835 27174 4881 27226
rect 4881 27174 4891 27226
rect 4915 27174 4945 27226
rect 4945 27174 4957 27226
rect 4957 27174 4971 27226
rect 4995 27174 5009 27226
rect 5009 27174 5021 27226
rect 5021 27174 5051 27226
rect 5075 27174 5085 27226
rect 5085 27174 5131 27226
rect 4835 27172 4891 27174
rect 4915 27172 4971 27174
rect 4995 27172 5051 27174
rect 5075 27172 5131 27174
rect 4175 26682 4231 26684
rect 4255 26682 4311 26684
rect 4335 26682 4391 26684
rect 4415 26682 4471 26684
rect 4175 26630 4221 26682
rect 4221 26630 4231 26682
rect 4255 26630 4285 26682
rect 4285 26630 4297 26682
rect 4297 26630 4311 26682
rect 4335 26630 4349 26682
rect 4349 26630 4361 26682
rect 4361 26630 4391 26682
rect 4415 26630 4425 26682
rect 4425 26630 4471 26682
rect 4175 26628 4231 26630
rect 4255 26628 4311 26630
rect 4335 26628 4391 26630
rect 4415 26628 4471 26630
rect 3422 25880 3478 25936
rect 1582 19896 1638 19952
rect 1582 19760 1638 19816
rect 938 19352 994 19408
rect 938 17176 994 17232
rect 1582 15952 1638 16008
rect 1398 15000 1454 15056
rect 1398 12824 1454 12880
rect 4835 26138 4891 26140
rect 4915 26138 4971 26140
rect 4995 26138 5051 26140
rect 5075 26138 5131 26140
rect 4835 26086 4881 26138
rect 4881 26086 4891 26138
rect 4915 26086 4945 26138
rect 4945 26086 4957 26138
rect 4957 26086 4971 26138
rect 4995 26086 5009 26138
rect 5009 26086 5021 26138
rect 5021 26086 5051 26138
rect 5075 26086 5085 26138
rect 5085 26086 5131 26138
rect 4835 26084 4891 26086
rect 4915 26084 4971 26086
rect 4995 26084 5051 26086
rect 5075 26084 5131 26086
rect 4175 25594 4231 25596
rect 4255 25594 4311 25596
rect 4335 25594 4391 25596
rect 4415 25594 4471 25596
rect 4175 25542 4221 25594
rect 4221 25542 4231 25594
rect 4255 25542 4285 25594
rect 4285 25542 4297 25594
rect 4297 25542 4311 25594
rect 4335 25542 4349 25594
rect 4349 25542 4361 25594
rect 4361 25542 4391 25594
rect 4415 25542 4425 25594
rect 4425 25542 4471 25594
rect 4175 25540 4231 25542
rect 4255 25540 4311 25542
rect 4335 25540 4391 25542
rect 4415 25540 4471 25542
rect 4175 24506 4231 24508
rect 4255 24506 4311 24508
rect 4335 24506 4391 24508
rect 4415 24506 4471 24508
rect 4175 24454 4221 24506
rect 4221 24454 4231 24506
rect 4255 24454 4285 24506
rect 4285 24454 4297 24506
rect 4297 24454 4311 24506
rect 4335 24454 4349 24506
rect 4349 24454 4361 24506
rect 4361 24454 4391 24506
rect 4415 24454 4425 24506
rect 4425 24454 4471 24506
rect 4175 24452 4231 24454
rect 4255 24452 4311 24454
rect 4335 24452 4391 24454
rect 4415 24452 4471 24454
rect 4835 25050 4891 25052
rect 4915 25050 4971 25052
rect 4995 25050 5051 25052
rect 5075 25050 5131 25052
rect 4835 24998 4881 25050
rect 4881 24998 4891 25050
rect 4915 24998 4945 25050
rect 4945 24998 4957 25050
rect 4957 24998 4971 25050
rect 4995 24998 5009 25050
rect 5009 24998 5021 25050
rect 5021 24998 5051 25050
rect 5075 24998 5085 25050
rect 5085 24998 5131 25050
rect 4835 24996 4891 24998
rect 4915 24996 4971 24998
rect 4995 24996 5051 24998
rect 5075 24996 5131 24998
rect 4835 23962 4891 23964
rect 4915 23962 4971 23964
rect 4995 23962 5051 23964
rect 5075 23962 5131 23964
rect 4835 23910 4881 23962
rect 4881 23910 4891 23962
rect 4915 23910 4945 23962
rect 4945 23910 4957 23962
rect 4957 23910 4971 23962
rect 4995 23910 5009 23962
rect 5009 23910 5021 23962
rect 5021 23910 5051 23962
rect 5075 23910 5085 23962
rect 5085 23910 5131 23962
rect 4835 23908 4891 23910
rect 4915 23908 4971 23910
rect 4995 23908 5051 23910
rect 5075 23908 5131 23910
rect 4175 23418 4231 23420
rect 4255 23418 4311 23420
rect 4335 23418 4391 23420
rect 4415 23418 4471 23420
rect 4175 23366 4221 23418
rect 4221 23366 4231 23418
rect 4255 23366 4285 23418
rect 4285 23366 4297 23418
rect 4297 23366 4311 23418
rect 4335 23366 4349 23418
rect 4349 23366 4361 23418
rect 4361 23366 4391 23418
rect 4415 23366 4425 23418
rect 4425 23366 4471 23418
rect 4175 23364 4231 23366
rect 4255 23364 4311 23366
rect 4335 23364 4391 23366
rect 4415 23364 4471 23366
rect 4175 22330 4231 22332
rect 4255 22330 4311 22332
rect 4335 22330 4391 22332
rect 4415 22330 4471 22332
rect 4175 22278 4221 22330
rect 4221 22278 4231 22330
rect 4255 22278 4285 22330
rect 4285 22278 4297 22330
rect 4297 22278 4311 22330
rect 4335 22278 4349 22330
rect 4349 22278 4361 22330
rect 4361 22278 4391 22330
rect 4415 22278 4425 22330
rect 4425 22278 4471 22330
rect 4175 22276 4231 22278
rect 4255 22276 4311 22278
rect 4335 22276 4391 22278
rect 4415 22276 4471 22278
rect 4835 22874 4891 22876
rect 4915 22874 4971 22876
rect 4995 22874 5051 22876
rect 5075 22874 5131 22876
rect 4835 22822 4881 22874
rect 4881 22822 4891 22874
rect 4915 22822 4945 22874
rect 4945 22822 4957 22874
rect 4957 22822 4971 22874
rect 4995 22822 5009 22874
rect 5009 22822 5021 22874
rect 5021 22822 5051 22874
rect 5075 22822 5085 22874
rect 5085 22822 5131 22874
rect 4835 22820 4891 22822
rect 4915 22820 4971 22822
rect 4995 22820 5051 22822
rect 5075 22820 5131 22822
rect 4066 21972 4068 21992
rect 4068 21972 4120 21992
rect 4120 21972 4122 21992
rect 4066 21936 4122 21972
rect 6182 23160 6238 23216
rect 4175 21242 4231 21244
rect 4255 21242 4311 21244
rect 4335 21242 4391 21244
rect 4415 21242 4471 21244
rect 4175 21190 4221 21242
rect 4221 21190 4231 21242
rect 4255 21190 4285 21242
rect 4285 21190 4297 21242
rect 4297 21190 4311 21242
rect 4335 21190 4349 21242
rect 4349 21190 4361 21242
rect 4361 21190 4391 21242
rect 4415 21190 4425 21242
rect 4425 21190 4471 21242
rect 4175 21188 4231 21190
rect 4255 21188 4311 21190
rect 4335 21188 4391 21190
rect 4415 21188 4471 21190
rect 5078 21972 5080 21992
rect 5080 21972 5132 21992
rect 5132 21972 5134 21992
rect 5078 21936 5134 21972
rect 4835 21786 4891 21788
rect 4915 21786 4971 21788
rect 4995 21786 5051 21788
rect 5075 21786 5131 21788
rect 4835 21734 4881 21786
rect 4881 21734 4891 21786
rect 4915 21734 4945 21786
rect 4945 21734 4957 21786
rect 4957 21734 4971 21786
rect 4995 21734 5009 21786
rect 5009 21734 5021 21786
rect 5021 21734 5051 21786
rect 5075 21734 5085 21786
rect 5085 21734 5131 21786
rect 4835 21732 4891 21734
rect 4915 21732 4971 21734
rect 4995 21732 5051 21734
rect 5075 21732 5131 21734
rect 4835 20698 4891 20700
rect 4915 20698 4971 20700
rect 4995 20698 5051 20700
rect 5075 20698 5131 20700
rect 4835 20646 4881 20698
rect 4881 20646 4891 20698
rect 4915 20646 4945 20698
rect 4945 20646 4957 20698
rect 4957 20646 4971 20698
rect 4995 20646 5009 20698
rect 5009 20646 5021 20698
rect 5021 20646 5051 20698
rect 5075 20646 5085 20698
rect 5085 20646 5131 20698
rect 4835 20644 4891 20646
rect 4915 20644 4971 20646
rect 4995 20644 5051 20646
rect 5075 20644 5131 20646
rect 4175 20154 4231 20156
rect 4255 20154 4311 20156
rect 4335 20154 4391 20156
rect 4415 20154 4471 20156
rect 4175 20102 4221 20154
rect 4221 20102 4231 20154
rect 4255 20102 4285 20154
rect 4285 20102 4297 20154
rect 4297 20102 4311 20154
rect 4335 20102 4349 20154
rect 4349 20102 4361 20154
rect 4361 20102 4391 20154
rect 4415 20102 4425 20154
rect 4425 20102 4471 20154
rect 4175 20100 4231 20102
rect 4255 20100 4311 20102
rect 4335 20100 4391 20102
rect 4415 20100 4471 20102
rect 4175 19066 4231 19068
rect 4255 19066 4311 19068
rect 4335 19066 4391 19068
rect 4415 19066 4471 19068
rect 4175 19014 4221 19066
rect 4221 19014 4231 19066
rect 4255 19014 4285 19066
rect 4285 19014 4297 19066
rect 4297 19014 4311 19066
rect 4335 19014 4349 19066
rect 4349 19014 4361 19066
rect 4361 19014 4391 19066
rect 4415 19014 4425 19066
rect 4425 19014 4471 19066
rect 4175 19012 4231 19014
rect 4255 19012 4311 19014
rect 4335 19012 4391 19014
rect 4415 19012 4471 19014
rect 4835 19610 4891 19612
rect 4915 19610 4971 19612
rect 4995 19610 5051 19612
rect 5075 19610 5131 19612
rect 4835 19558 4881 19610
rect 4881 19558 4891 19610
rect 4915 19558 4945 19610
rect 4945 19558 4957 19610
rect 4957 19558 4971 19610
rect 4995 19558 5009 19610
rect 5009 19558 5021 19610
rect 5021 19558 5051 19610
rect 5075 19558 5085 19610
rect 5085 19558 5131 19610
rect 4835 19556 4891 19558
rect 4915 19556 4971 19558
rect 4995 19556 5051 19558
rect 5075 19556 5131 19558
rect 9310 23740 9312 23760
rect 9312 23740 9364 23760
rect 9364 23740 9366 23760
rect 9310 23704 9366 23740
rect 9034 23296 9090 23352
rect 8942 23024 8998 23080
rect 9126 22616 9182 22672
rect 10322 23724 10378 23760
rect 10322 23704 10324 23724
rect 10324 23704 10376 23724
rect 10376 23704 10378 23724
rect 9770 23604 9772 23624
rect 9772 23604 9824 23624
rect 9824 23604 9826 23624
rect 9770 23568 9826 23604
rect 9862 23296 9918 23352
rect 9770 23060 9772 23080
rect 9772 23060 9824 23080
rect 9824 23060 9826 23080
rect 9770 23024 9826 23060
rect 5262 19352 5318 19408
rect 4835 18522 4891 18524
rect 4915 18522 4971 18524
rect 4995 18522 5051 18524
rect 5075 18522 5131 18524
rect 4835 18470 4881 18522
rect 4881 18470 4891 18522
rect 4915 18470 4945 18522
rect 4945 18470 4957 18522
rect 4957 18470 4971 18522
rect 4995 18470 5009 18522
rect 5009 18470 5021 18522
rect 5021 18470 5051 18522
rect 5075 18470 5085 18522
rect 5085 18470 5131 18522
rect 4835 18468 4891 18470
rect 4915 18468 4971 18470
rect 4995 18468 5051 18470
rect 5075 18468 5131 18470
rect 4175 17978 4231 17980
rect 4255 17978 4311 17980
rect 4335 17978 4391 17980
rect 4415 17978 4471 17980
rect 4175 17926 4221 17978
rect 4221 17926 4231 17978
rect 4255 17926 4285 17978
rect 4285 17926 4297 17978
rect 4297 17926 4311 17978
rect 4335 17926 4349 17978
rect 4349 17926 4361 17978
rect 4361 17926 4391 17978
rect 4415 17926 4425 17978
rect 4425 17926 4471 17978
rect 4175 17924 4231 17926
rect 4255 17924 4311 17926
rect 4335 17924 4391 17926
rect 4415 17924 4471 17926
rect 4835 17434 4891 17436
rect 4915 17434 4971 17436
rect 4995 17434 5051 17436
rect 5075 17434 5131 17436
rect 4835 17382 4881 17434
rect 4881 17382 4891 17434
rect 4915 17382 4945 17434
rect 4945 17382 4957 17434
rect 4957 17382 4971 17434
rect 4995 17382 5009 17434
rect 5009 17382 5021 17434
rect 5021 17382 5051 17434
rect 5075 17382 5085 17434
rect 5085 17382 5131 17434
rect 4835 17380 4891 17382
rect 4915 17380 4971 17382
rect 4995 17380 5051 17382
rect 5075 17380 5131 17382
rect 1398 10648 1454 10704
rect 938 8472 994 8528
rect 938 6316 994 6352
rect 938 6296 940 6316
rect 940 6296 992 6316
rect 992 6296 994 6316
rect 938 4120 994 4176
rect 938 1944 994 2000
rect 4175 16890 4231 16892
rect 4255 16890 4311 16892
rect 4335 16890 4391 16892
rect 4415 16890 4471 16892
rect 4175 16838 4221 16890
rect 4221 16838 4231 16890
rect 4255 16838 4285 16890
rect 4285 16838 4297 16890
rect 4297 16838 4311 16890
rect 4335 16838 4349 16890
rect 4349 16838 4361 16890
rect 4361 16838 4391 16890
rect 4415 16838 4425 16890
rect 4425 16838 4471 16890
rect 4175 16836 4231 16838
rect 4255 16836 4311 16838
rect 4335 16836 4391 16838
rect 4415 16836 4471 16838
rect 4835 16346 4891 16348
rect 4915 16346 4971 16348
rect 4995 16346 5051 16348
rect 5075 16346 5131 16348
rect 4835 16294 4881 16346
rect 4881 16294 4891 16346
rect 4915 16294 4945 16346
rect 4945 16294 4957 16346
rect 4957 16294 4971 16346
rect 4995 16294 5009 16346
rect 5009 16294 5021 16346
rect 5021 16294 5051 16346
rect 5075 16294 5085 16346
rect 5085 16294 5131 16346
rect 4835 16292 4891 16294
rect 4915 16292 4971 16294
rect 4995 16292 5051 16294
rect 5075 16292 5131 16294
rect 9678 22480 9734 22536
rect 9862 21956 9918 21992
rect 9862 21936 9864 21956
rect 9864 21936 9916 21956
rect 9916 21936 9918 21956
rect 11274 27226 11330 27228
rect 11354 27226 11410 27228
rect 11434 27226 11490 27228
rect 11514 27226 11570 27228
rect 11274 27174 11320 27226
rect 11320 27174 11330 27226
rect 11354 27174 11384 27226
rect 11384 27174 11396 27226
rect 11396 27174 11410 27226
rect 11434 27174 11448 27226
rect 11448 27174 11460 27226
rect 11460 27174 11490 27226
rect 11514 27174 11524 27226
rect 11524 27174 11570 27226
rect 11274 27172 11330 27174
rect 11354 27172 11410 27174
rect 11434 27172 11490 27174
rect 11514 27172 11570 27174
rect 10614 26682 10670 26684
rect 10694 26682 10750 26684
rect 10774 26682 10830 26684
rect 10854 26682 10910 26684
rect 10614 26630 10660 26682
rect 10660 26630 10670 26682
rect 10694 26630 10724 26682
rect 10724 26630 10736 26682
rect 10736 26630 10750 26682
rect 10774 26630 10788 26682
rect 10788 26630 10800 26682
rect 10800 26630 10830 26682
rect 10854 26630 10864 26682
rect 10864 26630 10910 26682
rect 10614 26628 10670 26630
rect 10694 26628 10750 26630
rect 10774 26628 10830 26630
rect 10854 26628 10910 26630
rect 10614 25594 10670 25596
rect 10694 25594 10750 25596
rect 10774 25594 10830 25596
rect 10854 25594 10910 25596
rect 10614 25542 10660 25594
rect 10660 25542 10670 25594
rect 10694 25542 10724 25594
rect 10724 25542 10736 25594
rect 10736 25542 10750 25594
rect 10774 25542 10788 25594
rect 10788 25542 10800 25594
rect 10800 25542 10830 25594
rect 10854 25542 10864 25594
rect 10864 25542 10910 25594
rect 10614 25540 10670 25542
rect 10694 25540 10750 25542
rect 10774 25540 10830 25542
rect 10854 25540 10910 25542
rect 11274 26138 11330 26140
rect 11354 26138 11410 26140
rect 11434 26138 11490 26140
rect 11514 26138 11570 26140
rect 11274 26086 11320 26138
rect 11320 26086 11330 26138
rect 11354 26086 11384 26138
rect 11384 26086 11396 26138
rect 11396 26086 11410 26138
rect 11434 26086 11448 26138
rect 11448 26086 11460 26138
rect 11460 26086 11490 26138
rect 11514 26086 11524 26138
rect 11524 26086 11570 26138
rect 11274 26084 11330 26086
rect 11354 26084 11410 26086
rect 11434 26084 11490 26086
rect 11514 26084 11570 26086
rect 11274 25050 11330 25052
rect 11354 25050 11410 25052
rect 11434 25050 11490 25052
rect 11514 25050 11570 25052
rect 11274 24998 11320 25050
rect 11320 24998 11330 25050
rect 11354 24998 11384 25050
rect 11384 24998 11396 25050
rect 11396 24998 11410 25050
rect 11434 24998 11448 25050
rect 11448 24998 11460 25050
rect 11460 24998 11490 25050
rect 11514 24998 11524 25050
rect 11524 24998 11570 25050
rect 11274 24996 11330 24998
rect 11354 24996 11410 24998
rect 11434 24996 11490 24998
rect 11514 24996 11570 24998
rect 10614 24506 10670 24508
rect 10694 24506 10750 24508
rect 10774 24506 10830 24508
rect 10854 24506 10910 24508
rect 10614 24454 10660 24506
rect 10660 24454 10670 24506
rect 10694 24454 10724 24506
rect 10724 24454 10736 24506
rect 10736 24454 10750 24506
rect 10774 24454 10788 24506
rect 10788 24454 10800 24506
rect 10800 24454 10830 24506
rect 10854 24454 10864 24506
rect 10864 24454 10910 24506
rect 10614 24452 10670 24454
rect 10694 24452 10750 24454
rect 10774 24452 10830 24454
rect 10854 24452 10910 24454
rect 10598 23604 10600 23624
rect 10600 23604 10652 23624
rect 10652 23604 10654 23624
rect 10598 23568 10654 23604
rect 10614 23418 10670 23420
rect 10694 23418 10750 23420
rect 10774 23418 10830 23420
rect 10854 23418 10910 23420
rect 10614 23366 10660 23418
rect 10660 23366 10670 23418
rect 10694 23366 10724 23418
rect 10724 23366 10736 23418
rect 10736 23366 10750 23418
rect 10774 23366 10788 23418
rect 10788 23366 10800 23418
rect 10800 23366 10830 23418
rect 10854 23366 10864 23418
rect 10864 23366 10910 23418
rect 10614 23364 10670 23366
rect 10694 23364 10750 23366
rect 10774 23364 10830 23366
rect 10854 23364 10910 23366
rect 4175 15802 4231 15804
rect 4255 15802 4311 15804
rect 4335 15802 4391 15804
rect 4415 15802 4471 15804
rect 4175 15750 4221 15802
rect 4221 15750 4231 15802
rect 4255 15750 4285 15802
rect 4285 15750 4297 15802
rect 4297 15750 4311 15802
rect 4335 15750 4349 15802
rect 4349 15750 4361 15802
rect 4361 15750 4391 15802
rect 4415 15750 4425 15802
rect 4425 15750 4471 15802
rect 4175 15748 4231 15750
rect 4255 15748 4311 15750
rect 4335 15748 4391 15750
rect 4415 15748 4471 15750
rect 4175 14714 4231 14716
rect 4255 14714 4311 14716
rect 4335 14714 4391 14716
rect 4415 14714 4471 14716
rect 4175 14662 4221 14714
rect 4221 14662 4231 14714
rect 4255 14662 4285 14714
rect 4285 14662 4297 14714
rect 4297 14662 4311 14714
rect 4335 14662 4349 14714
rect 4349 14662 4361 14714
rect 4361 14662 4391 14714
rect 4415 14662 4425 14714
rect 4425 14662 4471 14714
rect 4175 14660 4231 14662
rect 4255 14660 4311 14662
rect 4335 14660 4391 14662
rect 4415 14660 4471 14662
rect 4835 15258 4891 15260
rect 4915 15258 4971 15260
rect 4995 15258 5051 15260
rect 5075 15258 5131 15260
rect 4835 15206 4881 15258
rect 4881 15206 4891 15258
rect 4915 15206 4945 15258
rect 4945 15206 4957 15258
rect 4957 15206 4971 15258
rect 4995 15206 5009 15258
rect 5009 15206 5021 15258
rect 5021 15206 5051 15258
rect 5075 15206 5085 15258
rect 5085 15206 5131 15258
rect 4835 15204 4891 15206
rect 4915 15204 4971 15206
rect 4995 15204 5051 15206
rect 5075 15204 5131 15206
rect 4835 14170 4891 14172
rect 4915 14170 4971 14172
rect 4995 14170 5051 14172
rect 5075 14170 5131 14172
rect 4835 14118 4881 14170
rect 4881 14118 4891 14170
rect 4915 14118 4945 14170
rect 4945 14118 4957 14170
rect 4957 14118 4971 14170
rect 4995 14118 5009 14170
rect 5009 14118 5021 14170
rect 5021 14118 5051 14170
rect 5075 14118 5085 14170
rect 5085 14118 5131 14170
rect 4835 14116 4891 14118
rect 4915 14116 4971 14118
rect 4995 14116 5051 14118
rect 5075 14116 5131 14118
rect 7378 15952 7434 16008
rect 4175 13626 4231 13628
rect 4255 13626 4311 13628
rect 4335 13626 4391 13628
rect 4415 13626 4471 13628
rect 4175 13574 4221 13626
rect 4221 13574 4231 13626
rect 4255 13574 4285 13626
rect 4285 13574 4297 13626
rect 4297 13574 4311 13626
rect 4335 13574 4349 13626
rect 4349 13574 4361 13626
rect 4361 13574 4391 13626
rect 4415 13574 4425 13626
rect 4425 13574 4471 13626
rect 4175 13572 4231 13574
rect 4255 13572 4311 13574
rect 4335 13572 4391 13574
rect 4415 13572 4471 13574
rect 3974 12860 3976 12880
rect 3976 12860 4028 12880
rect 4028 12860 4030 12880
rect 3974 12824 4030 12860
rect 5078 13268 5080 13288
rect 5080 13268 5132 13288
rect 5132 13268 5134 13288
rect 5078 13232 5134 13268
rect 4835 13082 4891 13084
rect 4915 13082 4971 13084
rect 4995 13082 5051 13084
rect 5075 13082 5131 13084
rect 4835 13030 4881 13082
rect 4881 13030 4891 13082
rect 4915 13030 4945 13082
rect 4945 13030 4957 13082
rect 4957 13030 4971 13082
rect 4995 13030 5009 13082
rect 5009 13030 5021 13082
rect 5021 13030 5051 13082
rect 5075 13030 5085 13082
rect 5085 13030 5131 13082
rect 4835 13028 4891 13030
rect 4915 13028 4971 13030
rect 4995 13028 5051 13030
rect 5075 13028 5131 13030
rect 4175 12538 4231 12540
rect 4255 12538 4311 12540
rect 4335 12538 4391 12540
rect 4415 12538 4471 12540
rect 4175 12486 4221 12538
rect 4221 12486 4231 12538
rect 4255 12486 4285 12538
rect 4285 12486 4297 12538
rect 4297 12486 4311 12538
rect 4335 12486 4349 12538
rect 4349 12486 4361 12538
rect 4361 12486 4391 12538
rect 4415 12486 4425 12538
rect 4425 12486 4471 12538
rect 4175 12484 4231 12486
rect 4255 12484 4311 12486
rect 4335 12484 4391 12486
rect 4415 12484 4471 12486
rect 4835 11994 4891 11996
rect 4915 11994 4971 11996
rect 4995 11994 5051 11996
rect 5075 11994 5131 11996
rect 4835 11942 4881 11994
rect 4881 11942 4891 11994
rect 4915 11942 4945 11994
rect 4945 11942 4957 11994
rect 4957 11942 4971 11994
rect 4995 11942 5009 11994
rect 5009 11942 5021 11994
rect 5021 11942 5051 11994
rect 5075 11942 5085 11994
rect 5085 11942 5131 11994
rect 4835 11940 4891 11942
rect 4915 11940 4971 11942
rect 4995 11940 5051 11942
rect 5075 11940 5131 11942
rect 4175 11450 4231 11452
rect 4255 11450 4311 11452
rect 4335 11450 4391 11452
rect 4415 11450 4471 11452
rect 4175 11398 4221 11450
rect 4221 11398 4231 11450
rect 4255 11398 4285 11450
rect 4285 11398 4297 11450
rect 4297 11398 4311 11450
rect 4335 11398 4349 11450
rect 4349 11398 4361 11450
rect 4361 11398 4391 11450
rect 4415 11398 4425 11450
rect 4425 11398 4471 11450
rect 4175 11396 4231 11398
rect 4255 11396 4311 11398
rect 4335 11396 4391 11398
rect 4415 11396 4471 11398
rect 7654 13368 7710 13424
rect 8850 13268 8852 13288
rect 8852 13268 8904 13288
rect 8904 13268 8906 13288
rect 8850 13232 8906 13268
rect 9034 13232 9090 13288
rect 8850 12688 8906 12744
rect 10322 20032 10378 20088
rect 11274 23962 11330 23964
rect 11354 23962 11410 23964
rect 11434 23962 11490 23964
rect 11514 23962 11570 23964
rect 11274 23910 11320 23962
rect 11320 23910 11330 23962
rect 11354 23910 11384 23962
rect 11384 23910 11396 23962
rect 11396 23910 11410 23962
rect 11434 23910 11448 23962
rect 11448 23910 11460 23962
rect 11460 23910 11490 23962
rect 11514 23910 11524 23962
rect 11524 23910 11570 23962
rect 11274 23908 11330 23910
rect 11354 23908 11410 23910
rect 11434 23908 11490 23910
rect 11514 23908 11570 23910
rect 11426 23060 11428 23080
rect 11428 23060 11480 23080
rect 11480 23060 11482 23080
rect 10614 22330 10670 22332
rect 10694 22330 10750 22332
rect 10774 22330 10830 22332
rect 10854 22330 10910 22332
rect 10614 22278 10660 22330
rect 10660 22278 10670 22330
rect 10694 22278 10724 22330
rect 10724 22278 10736 22330
rect 10736 22278 10750 22330
rect 10774 22278 10788 22330
rect 10788 22278 10800 22330
rect 10800 22278 10830 22330
rect 10854 22278 10864 22330
rect 10864 22278 10910 22330
rect 10614 22276 10670 22278
rect 10694 22276 10750 22278
rect 10774 22276 10830 22278
rect 10854 22276 10910 22278
rect 11426 23024 11482 23060
rect 11274 22874 11330 22876
rect 11354 22874 11410 22876
rect 11434 22874 11490 22876
rect 11514 22874 11570 22876
rect 11274 22822 11320 22874
rect 11320 22822 11330 22874
rect 11354 22822 11384 22874
rect 11384 22822 11396 22874
rect 11396 22822 11410 22874
rect 11434 22822 11448 22874
rect 11448 22822 11460 22874
rect 11460 22822 11490 22874
rect 11514 22822 11524 22874
rect 11524 22822 11570 22874
rect 11274 22820 11330 22822
rect 11354 22820 11410 22822
rect 11434 22820 11490 22822
rect 11514 22820 11570 22822
rect 11058 22072 11114 22128
rect 11610 21972 11612 21992
rect 11612 21972 11664 21992
rect 11664 21972 11666 21992
rect 11610 21936 11666 21972
rect 10614 21242 10670 21244
rect 10694 21242 10750 21244
rect 10774 21242 10830 21244
rect 10854 21242 10910 21244
rect 10614 21190 10660 21242
rect 10660 21190 10670 21242
rect 10694 21190 10724 21242
rect 10724 21190 10736 21242
rect 10736 21190 10750 21242
rect 10774 21190 10788 21242
rect 10788 21190 10800 21242
rect 10800 21190 10830 21242
rect 10854 21190 10864 21242
rect 10864 21190 10910 21242
rect 10614 21188 10670 21190
rect 10694 21188 10750 21190
rect 10774 21188 10830 21190
rect 10854 21188 10910 21190
rect 11274 21786 11330 21788
rect 11354 21786 11410 21788
rect 11434 21786 11490 21788
rect 11514 21786 11570 21788
rect 11274 21734 11320 21786
rect 11320 21734 11330 21786
rect 11354 21734 11384 21786
rect 11384 21734 11396 21786
rect 11396 21734 11410 21786
rect 11434 21734 11448 21786
rect 11448 21734 11460 21786
rect 11460 21734 11490 21786
rect 11514 21734 11524 21786
rect 11524 21734 11570 21786
rect 11274 21732 11330 21734
rect 11354 21732 11410 21734
rect 11434 21732 11490 21734
rect 11514 21732 11570 21734
rect 11274 20698 11330 20700
rect 11354 20698 11410 20700
rect 11434 20698 11490 20700
rect 11514 20698 11570 20700
rect 11274 20646 11320 20698
rect 11320 20646 11330 20698
rect 11354 20646 11384 20698
rect 11384 20646 11396 20698
rect 11396 20646 11410 20698
rect 11434 20646 11448 20698
rect 11448 20646 11460 20698
rect 11460 20646 11490 20698
rect 11514 20646 11524 20698
rect 11524 20646 11570 20698
rect 11274 20644 11330 20646
rect 11354 20644 11410 20646
rect 11434 20644 11490 20646
rect 11514 20644 11570 20646
rect 11978 22616 12034 22672
rect 10414 19352 10470 19408
rect 10614 20154 10670 20156
rect 10694 20154 10750 20156
rect 10774 20154 10830 20156
rect 10854 20154 10910 20156
rect 10614 20102 10660 20154
rect 10660 20102 10670 20154
rect 10694 20102 10724 20154
rect 10724 20102 10736 20154
rect 10736 20102 10750 20154
rect 10774 20102 10788 20154
rect 10788 20102 10800 20154
rect 10800 20102 10830 20154
rect 10854 20102 10864 20154
rect 10864 20102 10910 20154
rect 10614 20100 10670 20102
rect 10694 20100 10750 20102
rect 10774 20100 10830 20102
rect 10854 20100 10910 20102
rect 10614 19066 10670 19068
rect 10694 19066 10750 19068
rect 10774 19066 10830 19068
rect 10854 19066 10910 19068
rect 10614 19014 10660 19066
rect 10660 19014 10670 19066
rect 10694 19014 10724 19066
rect 10724 19014 10736 19066
rect 10736 19014 10750 19066
rect 10774 19014 10788 19066
rect 10788 19014 10800 19066
rect 10800 19014 10830 19066
rect 10854 19014 10864 19066
rect 10864 19014 10910 19066
rect 10614 19012 10670 19014
rect 10694 19012 10750 19014
rect 10774 19012 10830 19014
rect 10854 19012 10910 19014
rect 9310 13232 9366 13288
rect 10614 17978 10670 17980
rect 10694 17978 10750 17980
rect 10774 17978 10830 17980
rect 10854 17978 10910 17980
rect 10614 17926 10660 17978
rect 10660 17926 10670 17978
rect 10694 17926 10724 17978
rect 10724 17926 10736 17978
rect 10736 17926 10750 17978
rect 10774 17926 10788 17978
rect 10788 17926 10800 17978
rect 10800 17926 10830 17978
rect 10854 17926 10864 17978
rect 10864 17926 10910 17978
rect 10614 17924 10670 17926
rect 10694 17924 10750 17926
rect 10774 17924 10830 17926
rect 10854 17924 10910 17926
rect 10614 16890 10670 16892
rect 10694 16890 10750 16892
rect 10774 16890 10830 16892
rect 10854 16890 10910 16892
rect 10614 16838 10660 16890
rect 10660 16838 10670 16890
rect 10694 16838 10724 16890
rect 10724 16838 10736 16890
rect 10736 16838 10750 16890
rect 10774 16838 10788 16890
rect 10788 16838 10800 16890
rect 10800 16838 10830 16890
rect 10854 16838 10864 16890
rect 10864 16838 10910 16890
rect 10614 16836 10670 16838
rect 10694 16836 10750 16838
rect 10774 16836 10830 16838
rect 10854 16836 10910 16838
rect 11794 19760 11850 19816
rect 11274 19610 11330 19612
rect 11354 19610 11410 19612
rect 11434 19610 11490 19612
rect 11514 19610 11570 19612
rect 11274 19558 11320 19610
rect 11320 19558 11330 19610
rect 11354 19558 11384 19610
rect 11384 19558 11396 19610
rect 11396 19558 11410 19610
rect 11434 19558 11448 19610
rect 11448 19558 11460 19610
rect 11460 19558 11490 19610
rect 11514 19558 11524 19610
rect 11524 19558 11570 19610
rect 11274 19556 11330 19558
rect 11354 19556 11410 19558
rect 11434 19556 11490 19558
rect 11514 19556 11570 19558
rect 11274 18522 11330 18524
rect 11354 18522 11410 18524
rect 11434 18522 11490 18524
rect 11514 18522 11570 18524
rect 11274 18470 11320 18522
rect 11320 18470 11330 18522
rect 11354 18470 11384 18522
rect 11384 18470 11396 18522
rect 11396 18470 11410 18522
rect 11434 18470 11448 18522
rect 11448 18470 11460 18522
rect 11460 18470 11490 18522
rect 11514 18470 11524 18522
rect 11524 18470 11570 18522
rect 11274 18468 11330 18470
rect 11354 18468 11410 18470
rect 11434 18468 11490 18470
rect 11514 18468 11570 18470
rect 11274 17434 11330 17436
rect 11354 17434 11410 17436
rect 11434 17434 11490 17436
rect 11514 17434 11570 17436
rect 11274 17382 11320 17434
rect 11320 17382 11330 17434
rect 11354 17382 11384 17434
rect 11384 17382 11396 17434
rect 11396 17382 11410 17434
rect 11434 17382 11448 17434
rect 11448 17382 11460 17434
rect 11460 17382 11490 17434
rect 11514 17382 11524 17434
rect 11524 17382 11570 17434
rect 11274 17380 11330 17382
rect 11354 17380 11410 17382
rect 11434 17380 11490 17382
rect 11514 17380 11570 17382
rect 11274 16346 11330 16348
rect 11354 16346 11410 16348
rect 11434 16346 11490 16348
rect 11514 16346 11570 16348
rect 11274 16294 11320 16346
rect 11320 16294 11330 16346
rect 11354 16294 11384 16346
rect 11384 16294 11396 16346
rect 11396 16294 11410 16346
rect 11434 16294 11448 16346
rect 11448 16294 11460 16346
rect 11460 16294 11490 16346
rect 11514 16294 11524 16346
rect 11524 16294 11570 16346
rect 11274 16292 11330 16294
rect 11354 16292 11410 16294
rect 11434 16292 11490 16294
rect 11514 16292 11570 16294
rect 11334 16108 11390 16144
rect 12714 22480 12770 22536
rect 15842 23160 15898 23216
rect 17713 27226 17769 27228
rect 17793 27226 17849 27228
rect 17873 27226 17929 27228
rect 17953 27226 18009 27228
rect 17713 27174 17759 27226
rect 17759 27174 17769 27226
rect 17793 27174 17823 27226
rect 17823 27174 17835 27226
rect 17835 27174 17849 27226
rect 17873 27174 17887 27226
rect 17887 27174 17899 27226
rect 17899 27174 17929 27226
rect 17953 27174 17963 27226
rect 17963 27174 18009 27226
rect 17713 27172 17769 27174
rect 17793 27172 17849 27174
rect 17873 27172 17929 27174
rect 17953 27172 18009 27174
rect 24152 27226 24208 27228
rect 24232 27226 24288 27228
rect 24312 27226 24368 27228
rect 24392 27226 24448 27228
rect 24152 27174 24198 27226
rect 24198 27174 24208 27226
rect 24232 27174 24262 27226
rect 24262 27174 24274 27226
rect 24274 27174 24288 27226
rect 24312 27174 24326 27226
rect 24326 27174 24338 27226
rect 24338 27174 24368 27226
rect 24392 27174 24402 27226
rect 24402 27174 24448 27226
rect 24152 27172 24208 27174
rect 24232 27172 24288 27174
rect 24312 27172 24368 27174
rect 24392 27172 24448 27174
rect 17053 26682 17109 26684
rect 17133 26682 17189 26684
rect 17213 26682 17269 26684
rect 17293 26682 17349 26684
rect 17053 26630 17099 26682
rect 17099 26630 17109 26682
rect 17133 26630 17163 26682
rect 17163 26630 17175 26682
rect 17175 26630 17189 26682
rect 17213 26630 17227 26682
rect 17227 26630 17239 26682
rect 17239 26630 17269 26682
rect 17293 26630 17303 26682
rect 17303 26630 17349 26682
rect 17053 26628 17109 26630
rect 17133 26628 17189 26630
rect 17213 26628 17269 26630
rect 17293 26628 17349 26630
rect 17713 26138 17769 26140
rect 17793 26138 17849 26140
rect 17873 26138 17929 26140
rect 17953 26138 18009 26140
rect 17713 26086 17759 26138
rect 17759 26086 17769 26138
rect 17793 26086 17823 26138
rect 17823 26086 17835 26138
rect 17835 26086 17849 26138
rect 17873 26086 17887 26138
rect 17887 26086 17899 26138
rect 17899 26086 17929 26138
rect 17953 26086 17963 26138
rect 17963 26086 18009 26138
rect 17713 26084 17769 26086
rect 17793 26084 17849 26086
rect 17873 26084 17929 26086
rect 17953 26084 18009 26086
rect 17053 25594 17109 25596
rect 17133 25594 17189 25596
rect 17213 25594 17269 25596
rect 17293 25594 17349 25596
rect 17053 25542 17099 25594
rect 17099 25542 17109 25594
rect 17133 25542 17163 25594
rect 17163 25542 17175 25594
rect 17175 25542 17189 25594
rect 17213 25542 17227 25594
rect 17227 25542 17239 25594
rect 17239 25542 17269 25594
rect 17293 25542 17303 25594
rect 17303 25542 17349 25594
rect 17053 25540 17109 25542
rect 17133 25540 17189 25542
rect 17213 25540 17269 25542
rect 17293 25540 17349 25542
rect 17713 25050 17769 25052
rect 17793 25050 17849 25052
rect 17873 25050 17929 25052
rect 17953 25050 18009 25052
rect 17713 24998 17759 25050
rect 17759 24998 17769 25050
rect 17793 24998 17823 25050
rect 17823 24998 17835 25050
rect 17835 24998 17849 25050
rect 17873 24998 17887 25050
rect 17887 24998 17899 25050
rect 17899 24998 17929 25050
rect 17953 24998 17963 25050
rect 17963 24998 18009 25050
rect 17713 24996 17769 24998
rect 17793 24996 17849 24998
rect 17873 24996 17929 24998
rect 17953 24996 18009 24998
rect 17053 24506 17109 24508
rect 17133 24506 17189 24508
rect 17213 24506 17269 24508
rect 17293 24506 17349 24508
rect 17053 24454 17099 24506
rect 17099 24454 17109 24506
rect 17133 24454 17163 24506
rect 17163 24454 17175 24506
rect 17175 24454 17189 24506
rect 17213 24454 17227 24506
rect 17227 24454 17239 24506
rect 17239 24454 17269 24506
rect 17293 24454 17303 24506
rect 17303 24454 17349 24506
rect 17053 24452 17109 24454
rect 17133 24452 17189 24454
rect 17213 24452 17269 24454
rect 17293 24452 17349 24454
rect 17713 23962 17769 23964
rect 17793 23962 17849 23964
rect 17873 23962 17929 23964
rect 17953 23962 18009 23964
rect 17713 23910 17759 23962
rect 17759 23910 17769 23962
rect 17793 23910 17823 23962
rect 17823 23910 17835 23962
rect 17835 23910 17849 23962
rect 17873 23910 17887 23962
rect 17887 23910 17899 23962
rect 17899 23910 17929 23962
rect 17953 23910 17963 23962
rect 17963 23910 18009 23962
rect 17713 23908 17769 23910
rect 17793 23908 17849 23910
rect 17873 23908 17929 23910
rect 17953 23908 18009 23910
rect 23492 26682 23548 26684
rect 23572 26682 23628 26684
rect 23652 26682 23708 26684
rect 23732 26682 23788 26684
rect 23492 26630 23538 26682
rect 23538 26630 23548 26682
rect 23572 26630 23602 26682
rect 23602 26630 23614 26682
rect 23614 26630 23628 26682
rect 23652 26630 23666 26682
rect 23666 26630 23678 26682
rect 23678 26630 23708 26682
rect 23732 26630 23742 26682
rect 23742 26630 23788 26682
rect 23492 26628 23548 26630
rect 23572 26628 23628 26630
rect 23652 26628 23708 26630
rect 23732 26628 23788 26630
rect 17053 23418 17109 23420
rect 17133 23418 17189 23420
rect 17213 23418 17269 23420
rect 17293 23418 17349 23420
rect 17053 23366 17099 23418
rect 17099 23366 17109 23418
rect 17133 23366 17163 23418
rect 17163 23366 17175 23418
rect 17175 23366 17189 23418
rect 17213 23366 17227 23418
rect 17227 23366 17239 23418
rect 17239 23366 17269 23418
rect 17293 23366 17303 23418
rect 17303 23366 17349 23418
rect 17053 23364 17109 23366
rect 17133 23364 17189 23366
rect 17213 23364 17269 23366
rect 17293 23364 17349 23366
rect 18234 23024 18290 23080
rect 17713 22874 17769 22876
rect 17793 22874 17849 22876
rect 17873 22874 17929 22876
rect 17953 22874 18009 22876
rect 17713 22822 17759 22874
rect 17759 22822 17769 22874
rect 17793 22822 17823 22874
rect 17823 22822 17835 22874
rect 17835 22822 17849 22874
rect 17873 22822 17887 22874
rect 17887 22822 17899 22874
rect 17899 22822 17929 22874
rect 17953 22822 17963 22874
rect 17963 22822 18009 22874
rect 17713 22820 17769 22822
rect 17793 22820 17849 22822
rect 17873 22820 17929 22822
rect 17953 22820 18009 22822
rect 14554 20712 14610 20768
rect 12254 19896 12310 19952
rect 11334 16088 11336 16108
rect 11336 16088 11388 16108
rect 11388 16088 11390 16108
rect 10614 15802 10670 15804
rect 10694 15802 10750 15804
rect 10774 15802 10830 15804
rect 10854 15802 10910 15804
rect 10614 15750 10660 15802
rect 10660 15750 10670 15802
rect 10694 15750 10724 15802
rect 10724 15750 10736 15802
rect 10736 15750 10750 15802
rect 10774 15750 10788 15802
rect 10788 15750 10800 15802
rect 10800 15750 10830 15802
rect 10854 15750 10864 15802
rect 10864 15750 10910 15802
rect 10614 15748 10670 15750
rect 10694 15748 10750 15750
rect 10774 15748 10830 15750
rect 10854 15748 10910 15750
rect 10614 14714 10670 14716
rect 10694 14714 10750 14716
rect 10774 14714 10830 14716
rect 10854 14714 10910 14716
rect 10614 14662 10660 14714
rect 10660 14662 10670 14714
rect 10694 14662 10724 14714
rect 10724 14662 10736 14714
rect 10736 14662 10750 14714
rect 10774 14662 10788 14714
rect 10788 14662 10800 14714
rect 10800 14662 10830 14714
rect 10854 14662 10864 14714
rect 10864 14662 10910 14714
rect 10614 14660 10670 14662
rect 10694 14660 10750 14662
rect 10774 14660 10830 14662
rect 10854 14660 10910 14662
rect 10614 13626 10670 13628
rect 10694 13626 10750 13628
rect 10774 13626 10830 13628
rect 10854 13626 10910 13628
rect 10614 13574 10660 13626
rect 10660 13574 10670 13626
rect 10694 13574 10724 13626
rect 10724 13574 10736 13626
rect 10736 13574 10750 13626
rect 10774 13574 10788 13626
rect 10788 13574 10800 13626
rect 10800 13574 10830 13626
rect 10854 13574 10864 13626
rect 10864 13574 10910 13626
rect 10614 13572 10670 13574
rect 10694 13572 10750 13574
rect 10774 13572 10830 13574
rect 10854 13572 10910 13574
rect 4066 11056 4122 11112
rect 4835 10906 4891 10908
rect 4915 10906 4971 10908
rect 4995 10906 5051 10908
rect 5075 10906 5131 10908
rect 4835 10854 4881 10906
rect 4881 10854 4891 10906
rect 4915 10854 4945 10906
rect 4945 10854 4957 10906
rect 4957 10854 4971 10906
rect 4995 10854 5009 10906
rect 5009 10854 5021 10906
rect 5021 10854 5051 10906
rect 5075 10854 5085 10906
rect 5085 10854 5131 10906
rect 4835 10852 4891 10854
rect 4915 10852 4971 10854
rect 4995 10852 5051 10854
rect 5075 10852 5131 10854
rect 4175 10362 4231 10364
rect 4255 10362 4311 10364
rect 4335 10362 4391 10364
rect 4415 10362 4471 10364
rect 4175 10310 4221 10362
rect 4221 10310 4231 10362
rect 4255 10310 4285 10362
rect 4285 10310 4297 10362
rect 4297 10310 4311 10362
rect 4335 10310 4349 10362
rect 4349 10310 4361 10362
rect 4361 10310 4391 10362
rect 4415 10310 4425 10362
rect 4425 10310 4471 10362
rect 4175 10308 4231 10310
rect 4255 10308 4311 10310
rect 4335 10308 4391 10310
rect 4415 10308 4471 10310
rect 4175 9274 4231 9276
rect 4255 9274 4311 9276
rect 4335 9274 4391 9276
rect 4415 9274 4471 9276
rect 4175 9222 4221 9274
rect 4221 9222 4231 9274
rect 4255 9222 4285 9274
rect 4285 9222 4297 9274
rect 4297 9222 4311 9274
rect 4335 9222 4349 9274
rect 4349 9222 4361 9274
rect 4361 9222 4391 9274
rect 4415 9222 4425 9274
rect 4425 9222 4471 9274
rect 4175 9220 4231 9222
rect 4255 9220 4311 9222
rect 4335 9220 4391 9222
rect 4415 9220 4471 9222
rect 4802 10004 4804 10024
rect 4804 10004 4856 10024
rect 4856 10004 4858 10024
rect 4802 9968 4858 10004
rect 4835 9818 4891 9820
rect 4915 9818 4971 9820
rect 4995 9818 5051 9820
rect 5075 9818 5131 9820
rect 4835 9766 4881 9818
rect 4881 9766 4891 9818
rect 4915 9766 4945 9818
rect 4945 9766 4957 9818
rect 4957 9766 4971 9818
rect 4995 9766 5009 9818
rect 5009 9766 5021 9818
rect 5021 9766 5051 9818
rect 5075 9766 5085 9818
rect 5085 9766 5131 9818
rect 4835 9764 4891 9766
rect 4915 9764 4971 9766
rect 4995 9764 5051 9766
rect 5075 9764 5131 9766
rect 5354 9968 5410 10024
rect 6734 11056 6790 11112
rect 4835 8730 4891 8732
rect 4915 8730 4971 8732
rect 4995 8730 5051 8732
rect 5075 8730 5131 8732
rect 4835 8678 4881 8730
rect 4881 8678 4891 8730
rect 4915 8678 4945 8730
rect 4945 8678 4957 8730
rect 4957 8678 4971 8730
rect 4995 8678 5009 8730
rect 5009 8678 5021 8730
rect 5021 8678 5051 8730
rect 5075 8678 5085 8730
rect 5085 8678 5131 8730
rect 4835 8676 4891 8678
rect 4915 8676 4971 8678
rect 4995 8676 5051 8678
rect 5075 8676 5131 8678
rect 4175 8186 4231 8188
rect 4255 8186 4311 8188
rect 4335 8186 4391 8188
rect 4415 8186 4471 8188
rect 4175 8134 4221 8186
rect 4221 8134 4231 8186
rect 4255 8134 4285 8186
rect 4285 8134 4297 8186
rect 4297 8134 4311 8186
rect 4335 8134 4349 8186
rect 4349 8134 4361 8186
rect 4361 8134 4391 8186
rect 4415 8134 4425 8186
rect 4425 8134 4471 8186
rect 4175 8132 4231 8134
rect 4255 8132 4311 8134
rect 4335 8132 4391 8134
rect 4415 8132 4471 8134
rect 4175 7098 4231 7100
rect 4255 7098 4311 7100
rect 4335 7098 4391 7100
rect 4415 7098 4471 7100
rect 4175 7046 4221 7098
rect 4221 7046 4231 7098
rect 4255 7046 4285 7098
rect 4285 7046 4297 7098
rect 4297 7046 4311 7098
rect 4335 7046 4349 7098
rect 4349 7046 4361 7098
rect 4361 7046 4391 7098
rect 4415 7046 4425 7098
rect 4425 7046 4471 7098
rect 4175 7044 4231 7046
rect 4255 7044 4311 7046
rect 4335 7044 4391 7046
rect 4415 7044 4471 7046
rect 4835 7642 4891 7644
rect 4915 7642 4971 7644
rect 4995 7642 5051 7644
rect 5075 7642 5131 7644
rect 4835 7590 4881 7642
rect 4881 7590 4891 7642
rect 4915 7590 4945 7642
rect 4945 7590 4957 7642
rect 4957 7590 4971 7642
rect 4995 7590 5009 7642
rect 5009 7590 5021 7642
rect 5021 7590 5051 7642
rect 5075 7590 5085 7642
rect 5085 7590 5131 7642
rect 4835 7588 4891 7590
rect 4915 7588 4971 7590
rect 4995 7588 5051 7590
rect 5075 7588 5131 7590
rect 4175 6010 4231 6012
rect 4255 6010 4311 6012
rect 4335 6010 4391 6012
rect 4415 6010 4471 6012
rect 4175 5958 4221 6010
rect 4221 5958 4231 6010
rect 4255 5958 4285 6010
rect 4285 5958 4297 6010
rect 4297 5958 4311 6010
rect 4335 5958 4349 6010
rect 4349 5958 4361 6010
rect 4361 5958 4391 6010
rect 4415 5958 4425 6010
rect 4425 5958 4471 6010
rect 4175 5956 4231 5958
rect 4255 5956 4311 5958
rect 4335 5956 4391 5958
rect 4415 5956 4471 5958
rect 4175 4922 4231 4924
rect 4255 4922 4311 4924
rect 4335 4922 4391 4924
rect 4415 4922 4471 4924
rect 4175 4870 4221 4922
rect 4221 4870 4231 4922
rect 4255 4870 4285 4922
rect 4285 4870 4297 4922
rect 4297 4870 4311 4922
rect 4335 4870 4349 4922
rect 4349 4870 4361 4922
rect 4361 4870 4391 4922
rect 4415 4870 4425 4922
rect 4425 4870 4471 4922
rect 4175 4868 4231 4870
rect 4255 4868 4311 4870
rect 4335 4868 4391 4870
rect 4415 4868 4471 4870
rect 4835 6554 4891 6556
rect 4915 6554 4971 6556
rect 4995 6554 5051 6556
rect 5075 6554 5131 6556
rect 4835 6502 4881 6554
rect 4881 6502 4891 6554
rect 4915 6502 4945 6554
rect 4945 6502 4957 6554
rect 4957 6502 4971 6554
rect 4995 6502 5009 6554
rect 5009 6502 5021 6554
rect 5021 6502 5051 6554
rect 5075 6502 5085 6554
rect 5085 6502 5131 6554
rect 4835 6500 4891 6502
rect 4915 6500 4971 6502
rect 4995 6500 5051 6502
rect 5075 6500 5131 6502
rect 4835 5466 4891 5468
rect 4915 5466 4971 5468
rect 4995 5466 5051 5468
rect 5075 5466 5131 5468
rect 4835 5414 4881 5466
rect 4881 5414 4891 5466
rect 4915 5414 4945 5466
rect 4945 5414 4957 5466
rect 4957 5414 4971 5466
rect 4995 5414 5009 5466
rect 5009 5414 5021 5466
rect 5021 5414 5051 5466
rect 5075 5414 5085 5466
rect 5085 5414 5131 5466
rect 4835 5412 4891 5414
rect 4915 5412 4971 5414
rect 4995 5412 5051 5414
rect 5075 5412 5131 5414
rect 4175 3834 4231 3836
rect 4255 3834 4311 3836
rect 4335 3834 4391 3836
rect 4415 3834 4471 3836
rect 4175 3782 4221 3834
rect 4221 3782 4231 3834
rect 4255 3782 4285 3834
rect 4285 3782 4297 3834
rect 4297 3782 4311 3834
rect 4335 3782 4349 3834
rect 4349 3782 4361 3834
rect 4361 3782 4391 3834
rect 4415 3782 4425 3834
rect 4425 3782 4471 3834
rect 4175 3780 4231 3782
rect 4255 3780 4311 3782
rect 4335 3780 4391 3782
rect 4415 3780 4471 3782
rect 4835 4378 4891 4380
rect 4915 4378 4971 4380
rect 4995 4378 5051 4380
rect 5075 4378 5131 4380
rect 4835 4326 4881 4378
rect 4881 4326 4891 4378
rect 4915 4326 4945 4378
rect 4945 4326 4957 4378
rect 4957 4326 4971 4378
rect 4995 4326 5009 4378
rect 5009 4326 5021 4378
rect 5021 4326 5051 4378
rect 5075 4326 5085 4378
rect 5085 4326 5131 4378
rect 4835 4324 4891 4326
rect 4915 4324 4971 4326
rect 4995 4324 5051 4326
rect 5075 4324 5131 4326
rect 4835 3290 4891 3292
rect 4915 3290 4971 3292
rect 4995 3290 5051 3292
rect 5075 3290 5131 3292
rect 4835 3238 4881 3290
rect 4881 3238 4891 3290
rect 4915 3238 4945 3290
rect 4945 3238 4957 3290
rect 4957 3238 4971 3290
rect 4995 3238 5009 3290
rect 5009 3238 5021 3290
rect 5021 3238 5051 3290
rect 5075 3238 5085 3290
rect 5085 3238 5131 3290
rect 4835 3236 4891 3238
rect 4915 3236 4971 3238
rect 4995 3236 5051 3238
rect 5075 3236 5131 3238
rect 10614 12538 10670 12540
rect 10694 12538 10750 12540
rect 10774 12538 10830 12540
rect 10854 12538 10910 12540
rect 10614 12486 10660 12538
rect 10660 12486 10670 12538
rect 10694 12486 10724 12538
rect 10724 12486 10736 12538
rect 10736 12486 10750 12538
rect 10774 12486 10788 12538
rect 10788 12486 10800 12538
rect 10800 12486 10830 12538
rect 10854 12486 10864 12538
rect 10864 12486 10910 12538
rect 10614 12484 10670 12486
rect 10694 12484 10750 12486
rect 10774 12484 10830 12486
rect 10854 12484 10910 12486
rect 11274 15258 11330 15260
rect 11354 15258 11410 15260
rect 11434 15258 11490 15260
rect 11514 15258 11570 15260
rect 11274 15206 11320 15258
rect 11320 15206 11330 15258
rect 11354 15206 11384 15258
rect 11384 15206 11396 15258
rect 11396 15206 11410 15258
rect 11434 15206 11448 15258
rect 11448 15206 11460 15258
rect 11460 15206 11490 15258
rect 11514 15206 11524 15258
rect 11524 15206 11570 15258
rect 11274 15204 11330 15206
rect 11354 15204 11410 15206
rect 11434 15204 11490 15206
rect 11514 15204 11570 15206
rect 11274 14170 11330 14172
rect 11354 14170 11410 14172
rect 11434 14170 11490 14172
rect 11514 14170 11570 14172
rect 11274 14118 11320 14170
rect 11320 14118 11330 14170
rect 11354 14118 11384 14170
rect 11384 14118 11396 14170
rect 11396 14118 11410 14170
rect 11434 14118 11448 14170
rect 11448 14118 11460 14170
rect 11460 14118 11490 14170
rect 11514 14118 11524 14170
rect 11524 14118 11570 14170
rect 11274 14116 11330 14118
rect 11354 14116 11410 14118
rect 11434 14116 11490 14118
rect 11514 14116 11570 14118
rect 11274 13082 11330 13084
rect 11354 13082 11410 13084
rect 11434 13082 11490 13084
rect 11514 13082 11570 13084
rect 11274 13030 11320 13082
rect 11320 13030 11330 13082
rect 11354 13030 11384 13082
rect 11384 13030 11396 13082
rect 11396 13030 11410 13082
rect 11434 13030 11448 13082
rect 11448 13030 11460 13082
rect 11460 13030 11490 13082
rect 11514 13030 11524 13082
rect 11524 13030 11570 13082
rect 11274 13028 11330 13030
rect 11354 13028 11410 13030
rect 11434 13028 11490 13030
rect 11514 13028 11570 13030
rect 9126 7248 9182 7304
rect 9586 6840 9642 6896
rect 8482 6740 8484 6760
rect 8484 6740 8536 6760
rect 8536 6740 8538 6760
rect 8482 6704 8538 6740
rect 8942 6316 8998 6352
rect 8942 6296 8944 6316
rect 8944 6296 8996 6316
rect 8996 6296 8998 6316
rect 9678 6568 9734 6624
rect 9954 6296 10010 6352
rect 10322 7248 10378 7304
rect 10230 6568 10286 6624
rect 13174 17176 13230 17232
rect 11274 11994 11330 11996
rect 11354 11994 11410 11996
rect 11434 11994 11490 11996
rect 11514 11994 11570 11996
rect 11274 11942 11320 11994
rect 11320 11942 11330 11994
rect 11354 11942 11384 11994
rect 11384 11942 11396 11994
rect 11396 11942 11410 11994
rect 11434 11942 11448 11994
rect 11448 11942 11460 11994
rect 11460 11942 11490 11994
rect 11514 11942 11524 11994
rect 11524 11942 11570 11994
rect 11274 11940 11330 11942
rect 11354 11940 11410 11942
rect 11434 11940 11490 11942
rect 11514 11940 11570 11942
rect 10614 11450 10670 11452
rect 10694 11450 10750 11452
rect 10774 11450 10830 11452
rect 10854 11450 10910 11452
rect 10614 11398 10660 11450
rect 10660 11398 10670 11450
rect 10694 11398 10724 11450
rect 10724 11398 10736 11450
rect 10736 11398 10750 11450
rect 10774 11398 10788 11450
rect 10788 11398 10800 11450
rect 10800 11398 10830 11450
rect 10854 11398 10864 11450
rect 10864 11398 10910 11450
rect 10614 11396 10670 11398
rect 10694 11396 10750 11398
rect 10774 11396 10830 11398
rect 10854 11396 10910 11398
rect 11274 10906 11330 10908
rect 11354 10906 11410 10908
rect 11434 10906 11490 10908
rect 11514 10906 11570 10908
rect 11274 10854 11320 10906
rect 11320 10854 11330 10906
rect 11354 10854 11384 10906
rect 11384 10854 11396 10906
rect 11396 10854 11410 10906
rect 11434 10854 11448 10906
rect 11448 10854 11460 10906
rect 11460 10854 11490 10906
rect 11514 10854 11524 10906
rect 11524 10854 11570 10906
rect 11274 10852 11330 10854
rect 11354 10852 11410 10854
rect 11434 10852 11490 10854
rect 11514 10852 11570 10854
rect 10614 10362 10670 10364
rect 10694 10362 10750 10364
rect 10774 10362 10830 10364
rect 10854 10362 10910 10364
rect 10614 10310 10660 10362
rect 10660 10310 10670 10362
rect 10694 10310 10724 10362
rect 10724 10310 10736 10362
rect 10736 10310 10750 10362
rect 10774 10310 10788 10362
rect 10788 10310 10800 10362
rect 10800 10310 10830 10362
rect 10854 10310 10864 10362
rect 10864 10310 10910 10362
rect 10614 10308 10670 10310
rect 10694 10308 10750 10310
rect 10774 10308 10830 10310
rect 10854 10308 10910 10310
rect 11274 9818 11330 9820
rect 11354 9818 11410 9820
rect 11434 9818 11490 9820
rect 11514 9818 11570 9820
rect 11274 9766 11320 9818
rect 11320 9766 11330 9818
rect 11354 9766 11384 9818
rect 11384 9766 11396 9818
rect 11396 9766 11410 9818
rect 11434 9766 11448 9818
rect 11448 9766 11460 9818
rect 11460 9766 11490 9818
rect 11514 9766 11524 9818
rect 11524 9766 11570 9818
rect 11274 9764 11330 9766
rect 11354 9764 11410 9766
rect 11434 9764 11490 9766
rect 11514 9764 11570 9766
rect 10614 9274 10670 9276
rect 10694 9274 10750 9276
rect 10774 9274 10830 9276
rect 10854 9274 10910 9276
rect 10614 9222 10660 9274
rect 10660 9222 10670 9274
rect 10694 9222 10724 9274
rect 10724 9222 10736 9274
rect 10736 9222 10750 9274
rect 10774 9222 10788 9274
rect 10788 9222 10800 9274
rect 10800 9222 10830 9274
rect 10854 9222 10864 9274
rect 10864 9222 10910 9274
rect 10614 9220 10670 9222
rect 10694 9220 10750 9222
rect 10774 9220 10830 9222
rect 10854 9220 10910 9222
rect 11058 9172 11114 9208
rect 11058 9152 11060 9172
rect 11060 9152 11112 9172
rect 11112 9152 11114 9172
rect 10782 8900 10838 8936
rect 10782 8880 10784 8900
rect 10784 8880 10836 8900
rect 10836 8880 10838 8900
rect 11274 8730 11330 8732
rect 11354 8730 11410 8732
rect 11434 8730 11490 8732
rect 11514 8730 11570 8732
rect 11274 8678 11320 8730
rect 11320 8678 11330 8730
rect 11354 8678 11384 8730
rect 11384 8678 11396 8730
rect 11396 8678 11410 8730
rect 11434 8678 11448 8730
rect 11448 8678 11460 8730
rect 11460 8678 11490 8730
rect 11514 8678 11524 8730
rect 11524 8678 11570 8730
rect 11274 8676 11330 8678
rect 11354 8676 11410 8678
rect 11434 8676 11490 8678
rect 11514 8676 11570 8678
rect 10614 8186 10670 8188
rect 10694 8186 10750 8188
rect 10774 8186 10830 8188
rect 10854 8186 10910 8188
rect 10614 8134 10660 8186
rect 10660 8134 10670 8186
rect 10694 8134 10724 8186
rect 10724 8134 10736 8186
rect 10736 8134 10750 8186
rect 10774 8134 10788 8186
rect 10788 8134 10800 8186
rect 10800 8134 10830 8186
rect 10854 8134 10864 8186
rect 10864 8134 10910 8186
rect 10614 8132 10670 8134
rect 10694 8132 10750 8134
rect 10774 8132 10830 8134
rect 10854 8132 10910 8134
rect 10598 7284 10600 7304
rect 10600 7284 10652 7304
rect 10652 7284 10654 7304
rect 10598 7248 10654 7284
rect 10614 7098 10670 7100
rect 10694 7098 10750 7100
rect 10774 7098 10830 7100
rect 10854 7098 10910 7100
rect 10614 7046 10660 7098
rect 10660 7046 10670 7098
rect 10694 7046 10724 7098
rect 10724 7046 10736 7098
rect 10736 7046 10750 7098
rect 10774 7046 10788 7098
rect 10788 7046 10800 7098
rect 10800 7046 10830 7098
rect 10854 7046 10864 7098
rect 10864 7046 10910 7098
rect 10614 7044 10670 7046
rect 10694 7044 10750 7046
rect 10774 7044 10830 7046
rect 10854 7044 10910 7046
rect 12530 13388 12586 13424
rect 12530 13368 12532 13388
rect 12532 13368 12584 13388
rect 12584 13368 12586 13388
rect 13174 16088 13230 16144
rect 13082 12824 13138 12880
rect 12990 9152 13046 9208
rect 11274 7642 11330 7644
rect 11354 7642 11410 7644
rect 11434 7642 11490 7644
rect 11514 7642 11570 7644
rect 11274 7590 11320 7642
rect 11320 7590 11330 7642
rect 11354 7590 11384 7642
rect 11384 7590 11396 7642
rect 11396 7590 11410 7642
rect 11434 7590 11448 7642
rect 11448 7590 11460 7642
rect 11460 7590 11490 7642
rect 11514 7590 11524 7642
rect 11524 7590 11570 7642
rect 11274 7588 11330 7590
rect 11354 7588 11410 7590
rect 11434 7588 11490 7590
rect 11514 7588 11570 7590
rect 11794 7404 11850 7440
rect 11794 7384 11796 7404
rect 11796 7384 11848 7404
rect 11848 7384 11850 7404
rect 10614 6010 10670 6012
rect 10694 6010 10750 6012
rect 10774 6010 10830 6012
rect 10854 6010 10910 6012
rect 10614 5958 10660 6010
rect 10660 5958 10670 6010
rect 10694 5958 10724 6010
rect 10724 5958 10736 6010
rect 10736 5958 10750 6010
rect 10774 5958 10788 6010
rect 10788 5958 10800 6010
rect 10800 5958 10830 6010
rect 10854 5958 10864 6010
rect 10864 5958 10910 6010
rect 10614 5956 10670 5958
rect 10694 5956 10750 5958
rect 10774 5956 10830 5958
rect 10854 5956 10910 5958
rect 4175 2746 4231 2748
rect 4255 2746 4311 2748
rect 4335 2746 4391 2748
rect 4415 2746 4471 2748
rect 4175 2694 4221 2746
rect 4221 2694 4231 2746
rect 4255 2694 4285 2746
rect 4285 2694 4297 2746
rect 4297 2694 4311 2746
rect 4335 2694 4349 2746
rect 4349 2694 4361 2746
rect 4361 2694 4391 2746
rect 4415 2694 4425 2746
rect 4425 2694 4471 2746
rect 4175 2692 4231 2694
rect 4255 2692 4311 2694
rect 4335 2692 4391 2694
rect 4415 2692 4471 2694
rect 10614 4922 10670 4924
rect 10694 4922 10750 4924
rect 10774 4922 10830 4924
rect 10854 4922 10910 4924
rect 10614 4870 10660 4922
rect 10660 4870 10670 4922
rect 10694 4870 10724 4922
rect 10724 4870 10736 4922
rect 10736 4870 10750 4922
rect 10774 4870 10788 4922
rect 10788 4870 10800 4922
rect 10800 4870 10830 4922
rect 10854 4870 10864 4922
rect 10864 4870 10910 4922
rect 10614 4868 10670 4870
rect 10694 4868 10750 4870
rect 10774 4868 10830 4870
rect 10854 4868 10910 4870
rect 11058 4528 11114 4584
rect 10614 3834 10670 3836
rect 10694 3834 10750 3836
rect 10774 3834 10830 3836
rect 10854 3834 10910 3836
rect 10614 3782 10660 3834
rect 10660 3782 10670 3834
rect 10694 3782 10724 3834
rect 10724 3782 10736 3834
rect 10736 3782 10750 3834
rect 10774 3782 10788 3834
rect 10788 3782 10800 3834
rect 10800 3782 10830 3834
rect 10854 3782 10864 3834
rect 10864 3782 10910 3834
rect 10614 3780 10670 3782
rect 10694 3780 10750 3782
rect 10774 3780 10830 3782
rect 10854 3780 10910 3782
rect 10614 2746 10670 2748
rect 10694 2746 10750 2748
rect 10774 2746 10830 2748
rect 10854 2746 10910 2748
rect 10614 2694 10660 2746
rect 10660 2694 10670 2746
rect 10694 2694 10724 2746
rect 10724 2694 10736 2746
rect 10736 2694 10750 2746
rect 10774 2694 10788 2746
rect 10788 2694 10800 2746
rect 10800 2694 10830 2746
rect 10854 2694 10864 2746
rect 10864 2694 10910 2746
rect 10614 2692 10670 2694
rect 10694 2692 10750 2694
rect 10774 2692 10830 2694
rect 10854 2692 10910 2694
rect 11274 6554 11330 6556
rect 11354 6554 11410 6556
rect 11434 6554 11490 6556
rect 11514 6554 11570 6556
rect 11274 6502 11320 6554
rect 11320 6502 11330 6554
rect 11354 6502 11384 6554
rect 11384 6502 11396 6554
rect 11396 6502 11410 6554
rect 11434 6502 11448 6554
rect 11448 6502 11460 6554
rect 11460 6502 11490 6554
rect 11514 6502 11524 6554
rect 11524 6502 11570 6554
rect 11274 6500 11330 6502
rect 11354 6500 11410 6502
rect 11434 6500 11490 6502
rect 11514 6500 11570 6502
rect 11274 5466 11330 5468
rect 11354 5466 11410 5468
rect 11434 5466 11490 5468
rect 11514 5466 11570 5468
rect 11274 5414 11320 5466
rect 11320 5414 11330 5466
rect 11354 5414 11384 5466
rect 11384 5414 11396 5466
rect 11396 5414 11410 5466
rect 11434 5414 11448 5466
rect 11448 5414 11460 5466
rect 11460 5414 11490 5466
rect 11514 5414 11524 5466
rect 11524 5414 11570 5466
rect 11274 5412 11330 5414
rect 11354 5412 11410 5414
rect 11434 5412 11490 5414
rect 11514 5412 11570 5414
rect 13266 8900 13322 8936
rect 13266 8880 13268 8900
rect 13268 8880 13320 8900
rect 13320 8880 13322 8900
rect 13634 5244 13636 5264
rect 13636 5244 13688 5264
rect 13688 5244 13690 5264
rect 13634 5208 13690 5244
rect 11274 4378 11330 4380
rect 11354 4378 11410 4380
rect 11434 4378 11490 4380
rect 11514 4378 11570 4380
rect 11274 4326 11320 4378
rect 11320 4326 11330 4378
rect 11354 4326 11384 4378
rect 11384 4326 11396 4378
rect 11396 4326 11410 4378
rect 11434 4326 11448 4378
rect 11448 4326 11460 4378
rect 11460 4326 11490 4378
rect 11514 4326 11524 4378
rect 11524 4326 11570 4378
rect 11274 4324 11330 4326
rect 11354 4324 11410 4326
rect 11434 4324 11490 4326
rect 11514 4324 11570 4326
rect 13082 4564 13084 4584
rect 13084 4564 13136 4584
rect 13136 4564 13138 4584
rect 13082 4528 13138 4564
rect 11274 3290 11330 3292
rect 11354 3290 11410 3292
rect 11434 3290 11490 3292
rect 11514 3290 11570 3292
rect 11274 3238 11320 3290
rect 11320 3238 11330 3290
rect 11354 3238 11384 3290
rect 11384 3238 11396 3290
rect 11396 3238 11410 3290
rect 11434 3238 11448 3290
rect 11448 3238 11460 3290
rect 11460 3238 11490 3290
rect 11514 3238 11524 3290
rect 11524 3238 11570 3290
rect 11274 3236 11330 3238
rect 11354 3236 11410 3238
rect 11434 3236 11490 3238
rect 11514 3236 11570 3238
rect 14462 12688 14518 12744
rect 15106 18808 15162 18864
rect 15474 17876 15530 17912
rect 15474 17856 15476 17876
rect 15476 17856 15528 17876
rect 15528 17856 15530 17876
rect 15842 20304 15898 20360
rect 16394 20324 16450 20360
rect 16394 20304 16396 20324
rect 16396 20304 16448 20324
rect 16448 20304 16450 20324
rect 15382 17332 15438 17368
rect 15382 17312 15384 17332
rect 15384 17312 15436 17332
rect 15436 17312 15438 17332
rect 15106 12724 15108 12744
rect 15108 12724 15160 12744
rect 15160 12724 15162 12744
rect 15106 12688 15162 12724
rect 15658 14340 15714 14376
rect 15658 14320 15660 14340
rect 15660 14320 15712 14340
rect 15712 14320 15714 14340
rect 15198 11736 15254 11792
rect 14370 6840 14426 6896
rect 14370 4392 14426 4448
rect 15198 6704 15254 6760
rect 15106 5228 15162 5264
rect 15106 5208 15108 5228
rect 15108 5208 15160 5228
rect 15160 5208 15162 5228
rect 17053 22330 17109 22332
rect 17133 22330 17189 22332
rect 17213 22330 17269 22332
rect 17293 22330 17349 22332
rect 17053 22278 17099 22330
rect 17099 22278 17109 22330
rect 17133 22278 17163 22330
rect 17163 22278 17175 22330
rect 17175 22278 17189 22330
rect 17213 22278 17227 22330
rect 17227 22278 17239 22330
rect 17239 22278 17269 22330
rect 17293 22278 17303 22330
rect 17303 22278 17349 22330
rect 17053 22276 17109 22278
rect 17133 22276 17189 22278
rect 17213 22276 17269 22278
rect 17293 22276 17349 22278
rect 18050 22072 18106 22128
rect 17713 21786 17769 21788
rect 17793 21786 17849 21788
rect 17873 21786 17929 21788
rect 17953 21786 18009 21788
rect 17713 21734 17759 21786
rect 17759 21734 17769 21786
rect 17793 21734 17823 21786
rect 17823 21734 17835 21786
rect 17835 21734 17849 21786
rect 17873 21734 17887 21786
rect 17887 21734 17899 21786
rect 17899 21734 17929 21786
rect 17953 21734 17963 21786
rect 17963 21734 18009 21786
rect 17713 21732 17769 21734
rect 17793 21732 17849 21734
rect 17873 21732 17929 21734
rect 17953 21732 18009 21734
rect 17053 21242 17109 21244
rect 17133 21242 17189 21244
rect 17213 21242 17269 21244
rect 17293 21242 17349 21244
rect 17053 21190 17099 21242
rect 17099 21190 17109 21242
rect 17133 21190 17163 21242
rect 17163 21190 17175 21242
rect 17175 21190 17189 21242
rect 17213 21190 17227 21242
rect 17227 21190 17239 21242
rect 17239 21190 17269 21242
rect 17293 21190 17303 21242
rect 17303 21190 17349 21242
rect 17053 21188 17109 21190
rect 17133 21188 17189 21190
rect 17213 21188 17269 21190
rect 17293 21188 17349 21190
rect 17038 20460 17094 20496
rect 17038 20440 17040 20460
rect 17040 20440 17092 20460
rect 17092 20440 17094 20460
rect 17053 20154 17109 20156
rect 17133 20154 17189 20156
rect 17213 20154 17269 20156
rect 17293 20154 17349 20156
rect 17053 20102 17099 20154
rect 17099 20102 17109 20154
rect 17133 20102 17163 20154
rect 17163 20102 17175 20154
rect 17175 20102 17189 20154
rect 17213 20102 17227 20154
rect 17227 20102 17239 20154
rect 17239 20102 17269 20154
rect 17293 20102 17303 20154
rect 17303 20102 17349 20154
rect 17053 20100 17109 20102
rect 17133 20100 17189 20102
rect 17213 20100 17269 20102
rect 17293 20100 17349 20102
rect 17053 19066 17109 19068
rect 17133 19066 17189 19068
rect 17213 19066 17269 19068
rect 17293 19066 17349 19068
rect 17053 19014 17099 19066
rect 17099 19014 17109 19066
rect 17133 19014 17163 19066
rect 17163 19014 17175 19066
rect 17175 19014 17189 19066
rect 17213 19014 17227 19066
rect 17227 19014 17239 19066
rect 17239 19014 17269 19066
rect 17293 19014 17303 19066
rect 17303 19014 17349 19066
rect 17053 19012 17109 19014
rect 17133 19012 17189 19014
rect 17213 19012 17269 19014
rect 17293 19012 17349 19014
rect 24152 26138 24208 26140
rect 24232 26138 24288 26140
rect 24312 26138 24368 26140
rect 24392 26138 24448 26140
rect 24152 26086 24198 26138
rect 24198 26086 24208 26138
rect 24232 26086 24262 26138
rect 24262 26086 24274 26138
rect 24274 26086 24288 26138
rect 24312 26086 24326 26138
rect 24326 26086 24338 26138
rect 24338 26086 24368 26138
rect 24392 26086 24402 26138
rect 24402 26086 24448 26138
rect 24152 26084 24208 26086
rect 24232 26084 24288 26086
rect 24312 26084 24368 26086
rect 24392 26084 24448 26086
rect 23492 25594 23548 25596
rect 23572 25594 23628 25596
rect 23652 25594 23708 25596
rect 23732 25594 23788 25596
rect 23492 25542 23538 25594
rect 23538 25542 23548 25594
rect 23572 25542 23602 25594
rect 23602 25542 23614 25594
rect 23614 25542 23628 25594
rect 23652 25542 23666 25594
rect 23666 25542 23678 25594
rect 23678 25542 23708 25594
rect 23732 25542 23742 25594
rect 23742 25542 23788 25594
rect 23492 25540 23548 25542
rect 23572 25540 23628 25542
rect 23652 25540 23708 25542
rect 23732 25540 23788 25542
rect 24152 25050 24208 25052
rect 24232 25050 24288 25052
rect 24312 25050 24368 25052
rect 24392 25050 24448 25052
rect 24152 24998 24198 25050
rect 24198 24998 24208 25050
rect 24232 24998 24262 25050
rect 24262 24998 24274 25050
rect 24274 24998 24288 25050
rect 24312 24998 24326 25050
rect 24326 24998 24338 25050
rect 24338 24998 24368 25050
rect 24392 24998 24402 25050
rect 24402 24998 24448 25050
rect 24152 24996 24208 24998
rect 24232 24996 24288 24998
rect 24312 24996 24368 24998
rect 24392 24996 24448 24998
rect 23492 24506 23548 24508
rect 23572 24506 23628 24508
rect 23652 24506 23708 24508
rect 23732 24506 23788 24508
rect 23492 24454 23538 24506
rect 23538 24454 23548 24506
rect 23572 24454 23602 24506
rect 23602 24454 23614 24506
rect 23614 24454 23628 24506
rect 23652 24454 23666 24506
rect 23666 24454 23678 24506
rect 23678 24454 23708 24506
rect 23732 24454 23742 24506
rect 23742 24454 23788 24506
rect 23492 24452 23548 24454
rect 23572 24452 23628 24454
rect 23652 24452 23708 24454
rect 23732 24452 23788 24454
rect 24152 23962 24208 23964
rect 24232 23962 24288 23964
rect 24312 23962 24368 23964
rect 24392 23962 24448 23964
rect 24152 23910 24198 23962
rect 24198 23910 24208 23962
rect 24232 23910 24262 23962
rect 24262 23910 24274 23962
rect 24274 23910 24288 23962
rect 24312 23910 24326 23962
rect 24326 23910 24338 23962
rect 24338 23910 24368 23962
rect 24392 23910 24402 23962
rect 24402 23910 24448 23962
rect 24152 23908 24208 23910
rect 24232 23908 24288 23910
rect 24312 23908 24368 23910
rect 24392 23908 24448 23910
rect 23492 23418 23548 23420
rect 23572 23418 23628 23420
rect 23652 23418 23708 23420
rect 23732 23418 23788 23420
rect 23492 23366 23538 23418
rect 23538 23366 23548 23418
rect 23572 23366 23602 23418
rect 23602 23366 23614 23418
rect 23614 23366 23628 23418
rect 23652 23366 23666 23418
rect 23666 23366 23678 23418
rect 23678 23366 23708 23418
rect 23732 23366 23742 23418
rect 23742 23366 23788 23418
rect 23492 23364 23548 23366
rect 23572 23364 23628 23366
rect 23652 23364 23708 23366
rect 23732 23364 23788 23366
rect 24152 22874 24208 22876
rect 24232 22874 24288 22876
rect 24312 22874 24368 22876
rect 24392 22874 24448 22876
rect 24152 22822 24198 22874
rect 24198 22822 24208 22874
rect 24232 22822 24262 22874
rect 24262 22822 24274 22874
rect 24274 22822 24288 22874
rect 24312 22822 24326 22874
rect 24326 22822 24338 22874
rect 24338 22822 24368 22874
rect 24392 22822 24402 22874
rect 24402 22822 24448 22874
rect 24152 22820 24208 22822
rect 24232 22820 24288 22822
rect 24312 22820 24368 22822
rect 24392 22820 24448 22822
rect 23492 22330 23548 22332
rect 23572 22330 23628 22332
rect 23652 22330 23708 22332
rect 23732 22330 23788 22332
rect 23492 22278 23538 22330
rect 23538 22278 23548 22330
rect 23572 22278 23602 22330
rect 23602 22278 23614 22330
rect 23614 22278 23628 22330
rect 23652 22278 23666 22330
rect 23666 22278 23678 22330
rect 23678 22278 23708 22330
rect 23732 22278 23742 22330
rect 23742 22278 23788 22330
rect 23492 22276 23548 22278
rect 23572 22276 23628 22278
rect 23652 22276 23708 22278
rect 23732 22276 23788 22278
rect 24152 21786 24208 21788
rect 24232 21786 24288 21788
rect 24312 21786 24368 21788
rect 24392 21786 24448 21788
rect 24152 21734 24198 21786
rect 24198 21734 24208 21786
rect 24232 21734 24262 21786
rect 24262 21734 24274 21786
rect 24274 21734 24288 21786
rect 24312 21734 24326 21786
rect 24326 21734 24338 21786
rect 24338 21734 24368 21786
rect 24392 21734 24402 21786
rect 24402 21734 24448 21786
rect 24152 21732 24208 21734
rect 24232 21732 24288 21734
rect 24312 21732 24368 21734
rect 24392 21732 24448 21734
rect 23492 21242 23548 21244
rect 23572 21242 23628 21244
rect 23652 21242 23708 21244
rect 23732 21242 23788 21244
rect 23492 21190 23538 21242
rect 23538 21190 23548 21242
rect 23572 21190 23602 21242
rect 23602 21190 23614 21242
rect 23614 21190 23628 21242
rect 23652 21190 23666 21242
rect 23666 21190 23678 21242
rect 23678 21190 23708 21242
rect 23732 21190 23742 21242
rect 23742 21190 23788 21242
rect 23492 21188 23548 21190
rect 23572 21188 23628 21190
rect 23652 21188 23708 21190
rect 23732 21188 23788 21190
rect 17713 20698 17769 20700
rect 17793 20698 17849 20700
rect 17873 20698 17929 20700
rect 17953 20698 18009 20700
rect 17713 20646 17759 20698
rect 17759 20646 17769 20698
rect 17793 20646 17823 20698
rect 17823 20646 17835 20698
rect 17835 20646 17849 20698
rect 17873 20646 17887 20698
rect 17887 20646 17899 20698
rect 17899 20646 17929 20698
rect 17953 20646 17963 20698
rect 17963 20646 18009 20698
rect 17713 20644 17769 20646
rect 17793 20644 17849 20646
rect 17873 20644 17929 20646
rect 17953 20644 18009 20646
rect 24152 20698 24208 20700
rect 24232 20698 24288 20700
rect 24312 20698 24368 20700
rect 24392 20698 24448 20700
rect 24152 20646 24198 20698
rect 24198 20646 24208 20698
rect 24232 20646 24262 20698
rect 24262 20646 24274 20698
rect 24274 20646 24288 20698
rect 24312 20646 24326 20698
rect 24326 20646 24338 20698
rect 24338 20646 24368 20698
rect 24392 20646 24402 20698
rect 24402 20646 24448 20698
rect 24152 20644 24208 20646
rect 24232 20644 24288 20646
rect 24312 20644 24368 20646
rect 24392 20644 24448 20646
rect 16118 4004 16174 4040
rect 16118 3984 16120 4004
rect 16120 3984 16172 4004
rect 16172 3984 16174 4004
rect 17053 17978 17109 17980
rect 17133 17978 17189 17980
rect 17213 17978 17269 17980
rect 17293 17978 17349 17980
rect 17053 17926 17099 17978
rect 17099 17926 17109 17978
rect 17133 17926 17163 17978
rect 17163 17926 17175 17978
rect 17175 17926 17189 17978
rect 17213 17926 17227 17978
rect 17227 17926 17239 17978
rect 17239 17926 17269 17978
rect 17293 17926 17303 17978
rect 17303 17926 17349 17978
rect 17053 17924 17109 17926
rect 17133 17924 17189 17926
rect 17213 17924 17269 17926
rect 17293 17924 17349 17926
rect 17053 16890 17109 16892
rect 17133 16890 17189 16892
rect 17213 16890 17269 16892
rect 17293 16890 17349 16892
rect 17053 16838 17099 16890
rect 17099 16838 17109 16890
rect 17133 16838 17163 16890
rect 17163 16838 17175 16890
rect 17175 16838 17189 16890
rect 17213 16838 17227 16890
rect 17227 16838 17239 16890
rect 17239 16838 17269 16890
rect 17293 16838 17303 16890
rect 17303 16838 17349 16890
rect 17053 16836 17109 16838
rect 17133 16836 17189 16838
rect 17213 16836 17269 16838
rect 17293 16836 17349 16838
rect 17406 16088 17462 16144
rect 17053 15802 17109 15804
rect 17133 15802 17189 15804
rect 17213 15802 17269 15804
rect 17293 15802 17349 15804
rect 17053 15750 17099 15802
rect 17099 15750 17109 15802
rect 17133 15750 17163 15802
rect 17163 15750 17175 15802
rect 17175 15750 17189 15802
rect 17213 15750 17227 15802
rect 17227 15750 17239 15802
rect 17239 15750 17269 15802
rect 17293 15750 17303 15802
rect 17303 15750 17349 15802
rect 17053 15748 17109 15750
rect 17133 15748 17189 15750
rect 17213 15748 17269 15750
rect 17293 15748 17349 15750
rect 17053 14714 17109 14716
rect 17133 14714 17189 14716
rect 17213 14714 17269 14716
rect 17293 14714 17349 14716
rect 17053 14662 17099 14714
rect 17099 14662 17109 14714
rect 17133 14662 17163 14714
rect 17163 14662 17175 14714
rect 17175 14662 17189 14714
rect 17213 14662 17227 14714
rect 17227 14662 17239 14714
rect 17239 14662 17269 14714
rect 17293 14662 17303 14714
rect 17303 14662 17349 14714
rect 17053 14660 17109 14662
rect 17133 14660 17189 14662
rect 17213 14660 17269 14662
rect 17293 14660 17349 14662
rect 17222 14456 17278 14512
rect 17713 19610 17769 19612
rect 17793 19610 17849 19612
rect 17873 19610 17929 19612
rect 17953 19610 18009 19612
rect 17713 19558 17759 19610
rect 17759 19558 17769 19610
rect 17793 19558 17823 19610
rect 17823 19558 17835 19610
rect 17835 19558 17849 19610
rect 17873 19558 17887 19610
rect 17887 19558 17899 19610
rect 17899 19558 17929 19610
rect 17953 19558 17963 19610
rect 17963 19558 18009 19610
rect 17713 19556 17769 19558
rect 17793 19556 17849 19558
rect 17873 19556 17929 19558
rect 17953 19556 18009 19558
rect 17958 18808 18014 18864
rect 17713 18522 17769 18524
rect 17793 18522 17849 18524
rect 17873 18522 17929 18524
rect 17953 18522 18009 18524
rect 17713 18470 17759 18522
rect 17759 18470 17769 18522
rect 17793 18470 17823 18522
rect 17823 18470 17835 18522
rect 17835 18470 17849 18522
rect 17873 18470 17887 18522
rect 17887 18470 17899 18522
rect 17899 18470 17929 18522
rect 17953 18470 17963 18522
rect 17963 18470 18009 18522
rect 17713 18468 17769 18470
rect 17793 18468 17849 18470
rect 17873 18468 17929 18470
rect 17953 18468 18009 18470
rect 17713 17434 17769 17436
rect 17793 17434 17849 17436
rect 17873 17434 17929 17436
rect 17953 17434 18009 17436
rect 17713 17382 17759 17434
rect 17759 17382 17769 17434
rect 17793 17382 17823 17434
rect 17823 17382 17835 17434
rect 17835 17382 17849 17434
rect 17873 17382 17887 17434
rect 17887 17382 17899 17434
rect 17899 17382 17929 17434
rect 17953 17382 17963 17434
rect 17963 17382 18009 17434
rect 17713 17380 17769 17382
rect 17793 17380 17849 17382
rect 17873 17380 17929 17382
rect 17953 17380 18009 17382
rect 17713 16346 17769 16348
rect 17793 16346 17849 16348
rect 17873 16346 17929 16348
rect 17953 16346 18009 16348
rect 17713 16294 17759 16346
rect 17759 16294 17769 16346
rect 17793 16294 17823 16346
rect 17823 16294 17835 16346
rect 17835 16294 17849 16346
rect 17873 16294 17887 16346
rect 17887 16294 17899 16346
rect 17899 16294 17929 16346
rect 17953 16294 17963 16346
rect 17963 16294 18009 16346
rect 17713 16292 17769 16294
rect 17793 16292 17849 16294
rect 17873 16292 17929 16294
rect 17953 16292 18009 16294
rect 17682 16088 17738 16144
rect 26146 25880 26202 25936
rect 25502 20304 25558 20360
rect 23492 20154 23548 20156
rect 23572 20154 23628 20156
rect 23652 20154 23708 20156
rect 23732 20154 23788 20156
rect 23492 20102 23538 20154
rect 23538 20102 23548 20154
rect 23572 20102 23602 20154
rect 23602 20102 23614 20154
rect 23614 20102 23628 20154
rect 23652 20102 23666 20154
rect 23666 20102 23678 20154
rect 23678 20102 23708 20154
rect 23732 20102 23742 20154
rect 23742 20102 23788 20154
rect 23492 20100 23548 20102
rect 23572 20100 23628 20102
rect 23652 20100 23708 20102
rect 23732 20100 23788 20102
rect 18786 17176 18842 17232
rect 18418 16108 18474 16144
rect 18418 16088 18420 16108
rect 18420 16088 18472 16108
rect 18472 16088 18474 16108
rect 17713 15258 17769 15260
rect 17793 15258 17849 15260
rect 17873 15258 17929 15260
rect 17953 15258 18009 15260
rect 17713 15206 17759 15258
rect 17759 15206 17769 15258
rect 17793 15206 17823 15258
rect 17823 15206 17835 15258
rect 17835 15206 17849 15258
rect 17873 15206 17887 15258
rect 17887 15206 17899 15258
rect 17899 15206 17929 15258
rect 17953 15206 17963 15258
rect 17963 15206 18009 15258
rect 17713 15204 17769 15206
rect 17793 15204 17849 15206
rect 17873 15204 17929 15206
rect 17953 15204 18009 15206
rect 17053 13626 17109 13628
rect 17133 13626 17189 13628
rect 17213 13626 17269 13628
rect 17293 13626 17349 13628
rect 17053 13574 17099 13626
rect 17099 13574 17109 13626
rect 17133 13574 17163 13626
rect 17163 13574 17175 13626
rect 17175 13574 17189 13626
rect 17213 13574 17227 13626
rect 17227 13574 17239 13626
rect 17239 13574 17269 13626
rect 17293 13574 17303 13626
rect 17303 13574 17349 13626
rect 17053 13572 17109 13574
rect 17133 13572 17189 13574
rect 17213 13572 17269 13574
rect 17293 13572 17349 13574
rect 17053 12538 17109 12540
rect 17133 12538 17189 12540
rect 17213 12538 17269 12540
rect 17293 12538 17349 12540
rect 17053 12486 17099 12538
rect 17099 12486 17109 12538
rect 17133 12486 17163 12538
rect 17163 12486 17175 12538
rect 17175 12486 17189 12538
rect 17213 12486 17227 12538
rect 17227 12486 17239 12538
rect 17239 12486 17269 12538
rect 17293 12486 17303 12538
rect 17303 12486 17349 12538
rect 17053 12484 17109 12486
rect 17133 12484 17189 12486
rect 17213 12484 17269 12486
rect 17293 12484 17349 12486
rect 17958 14456 18014 14512
rect 17713 14170 17769 14172
rect 17793 14170 17849 14172
rect 17873 14170 17929 14172
rect 17953 14170 18009 14172
rect 17713 14118 17759 14170
rect 17759 14118 17769 14170
rect 17793 14118 17823 14170
rect 17823 14118 17835 14170
rect 17835 14118 17849 14170
rect 17873 14118 17887 14170
rect 17887 14118 17899 14170
rect 17899 14118 17929 14170
rect 17953 14118 17963 14170
rect 17963 14118 18009 14170
rect 17713 14116 17769 14118
rect 17793 14116 17849 14118
rect 17873 14116 17929 14118
rect 17953 14116 18009 14118
rect 18326 14456 18382 14512
rect 18786 14320 18842 14376
rect 19062 14492 19064 14512
rect 19064 14492 19116 14512
rect 19116 14492 19118 14512
rect 19062 14456 19118 14492
rect 17713 13082 17769 13084
rect 17793 13082 17849 13084
rect 17873 13082 17929 13084
rect 17953 13082 18009 13084
rect 17713 13030 17759 13082
rect 17759 13030 17769 13082
rect 17793 13030 17823 13082
rect 17823 13030 17835 13082
rect 17835 13030 17849 13082
rect 17873 13030 17887 13082
rect 17887 13030 17899 13082
rect 17899 13030 17929 13082
rect 17953 13030 17963 13082
rect 17963 13030 18009 13082
rect 17713 13028 17769 13030
rect 17793 13028 17849 13030
rect 17873 13028 17929 13030
rect 17953 13028 18009 13030
rect 24152 19610 24208 19612
rect 24232 19610 24288 19612
rect 24312 19610 24368 19612
rect 24392 19610 24448 19612
rect 24152 19558 24198 19610
rect 24198 19558 24208 19610
rect 24232 19558 24262 19610
rect 24262 19558 24274 19610
rect 24274 19558 24288 19610
rect 24312 19558 24326 19610
rect 24326 19558 24338 19610
rect 24338 19558 24368 19610
rect 24392 19558 24402 19610
rect 24402 19558 24448 19610
rect 24152 19556 24208 19558
rect 24232 19556 24288 19558
rect 24312 19556 24368 19558
rect 24392 19556 24448 19558
rect 23492 19066 23548 19068
rect 23572 19066 23628 19068
rect 23652 19066 23708 19068
rect 23732 19066 23788 19068
rect 23492 19014 23538 19066
rect 23538 19014 23548 19066
rect 23572 19014 23602 19066
rect 23602 19014 23614 19066
rect 23614 19014 23628 19066
rect 23652 19014 23666 19066
rect 23666 19014 23678 19066
rect 23678 19014 23708 19066
rect 23732 19014 23742 19066
rect 23742 19014 23788 19066
rect 23492 19012 23548 19014
rect 23572 19012 23628 19014
rect 23652 19012 23708 19014
rect 23732 19012 23788 19014
rect 26514 18536 26570 18592
rect 24152 18522 24208 18524
rect 24232 18522 24288 18524
rect 24312 18522 24368 18524
rect 24392 18522 24448 18524
rect 24152 18470 24198 18522
rect 24198 18470 24208 18522
rect 24232 18470 24262 18522
rect 24262 18470 24274 18522
rect 24274 18470 24288 18522
rect 24312 18470 24326 18522
rect 24326 18470 24338 18522
rect 24338 18470 24368 18522
rect 24392 18470 24402 18522
rect 24402 18470 24448 18522
rect 24152 18468 24208 18470
rect 24232 18468 24288 18470
rect 24312 18468 24368 18470
rect 24392 18468 24448 18470
rect 23492 17978 23548 17980
rect 23572 17978 23628 17980
rect 23652 17978 23708 17980
rect 23732 17978 23788 17980
rect 23492 17926 23538 17978
rect 23538 17926 23548 17978
rect 23572 17926 23602 17978
rect 23602 17926 23614 17978
rect 23614 17926 23628 17978
rect 23652 17926 23666 17978
rect 23666 17926 23678 17978
rect 23678 17926 23708 17978
rect 23732 17926 23742 17978
rect 23742 17926 23788 17978
rect 23492 17924 23548 17926
rect 23572 17924 23628 17926
rect 23652 17924 23708 17926
rect 23732 17924 23788 17926
rect 16854 11756 16910 11792
rect 17713 11994 17769 11996
rect 17793 11994 17849 11996
rect 17873 11994 17929 11996
rect 17953 11994 18009 11996
rect 17713 11942 17759 11994
rect 17759 11942 17769 11994
rect 17793 11942 17823 11994
rect 17823 11942 17835 11994
rect 17835 11942 17849 11994
rect 17873 11942 17887 11994
rect 17887 11942 17899 11994
rect 17899 11942 17929 11994
rect 17953 11942 17963 11994
rect 17963 11942 18009 11994
rect 17713 11940 17769 11942
rect 17793 11940 17849 11942
rect 17873 11940 17929 11942
rect 17953 11940 18009 11942
rect 16854 11736 16856 11756
rect 16856 11736 16908 11756
rect 16908 11736 16910 11756
rect 17053 11450 17109 11452
rect 17133 11450 17189 11452
rect 17213 11450 17269 11452
rect 17293 11450 17349 11452
rect 17053 11398 17099 11450
rect 17099 11398 17109 11450
rect 17133 11398 17163 11450
rect 17163 11398 17175 11450
rect 17175 11398 17189 11450
rect 17213 11398 17227 11450
rect 17227 11398 17239 11450
rect 17239 11398 17269 11450
rect 17293 11398 17303 11450
rect 17303 11398 17349 11450
rect 17053 11396 17109 11398
rect 17133 11396 17189 11398
rect 17213 11396 17269 11398
rect 17293 11396 17349 11398
rect 24152 17434 24208 17436
rect 24232 17434 24288 17436
rect 24312 17434 24368 17436
rect 24392 17434 24448 17436
rect 24152 17382 24198 17434
rect 24198 17382 24208 17434
rect 24232 17382 24262 17434
rect 24262 17382 24274 17434
rect 24274 17382 24288 17434
rect 24312 17382 24326 17434
rect 24326 17382 24338 17434
rect 24338 17382 24368 17434
rect 24392 17382 24402 17434
rect 24402 17382 24448 17434
rect 24152 17380 24208 17382
rect 24232 17380 24288 17382
rect 24312 17380 24368 17382
rect 24392 17380 24448 17382
rect 23492 16890 23548 16892
rect 23572 16890 23628 16892
rect 23652 16890 23708 16892
rect 23732 16890 23788 16892
rect 23492 16838 23538 16890
rect 23538 16838 23548 16890
rect 23572 16838 23602 16890
rect 23602 16838 23614 16890
rect 23614 16838 23628 16890
rect 23652 16838 23666 16890
rect 23666 16838 23678 16890
rect 23678 16838 23708 16890
rect 23732 16838 23742 16890
rect 23742 16838 23788 16890
rect 23492 16836 23548 16838
rect 23572 16836 23628 16838
rect 23652 16836 23708 16838
rect 23732 16836 23788 16838
rect 20994 13232 21050 13288
rect 18786 11736 18842 11792
rect 17713 10906 17769 10908
rect 17793 10906 17849 10908
rect 17873 10906 17929 10908
rect 17953 10906 18009 10908
rect 17713 10854 17759 10906
rect 17759 10854 17769 10906
rect 17793 10854 17823 10906
rect 17823 10854 17835 10906
rect 17835 10854 17849 10906
rect 17873 10854 17887 10906
rect 17887 10854 17899 10906
rect 17899 10854 17929 10906
rect 17953 10854 17963 10906
rect 17963 10854 18009 10906
rect 17713 10852 17769 10854
rect 17793 10852 17849 10854
rect 17873 10852 17929 10854
rect 17953 10852 18009 10854
rect 23492 15802 23548 15804
rect 23572 15802 23628 15804
rect 23652 15802 23708 15804
rect 23732 15802 23788 15804
rect 23492 15750 23538 15802
rect 23538 15750 23548 15802
rect 23572 15750 23602 15802
rect 23602 15750 23614 15802
rect 23614 15750 23628 15802
rect 23652 15750 23666 15802
rect 23666 15750 23678 15802
rect 23678 15750 23708 15802
rect 23732 15750 23742 15802
rect 23742 15750 23788 15802
rect 23492 15748 23548 15750
rect 23572 15748 23628 15750
rect 23652 15748 23708 15750
rect 23732 15748 23788 15750
rect 24152 16346 24208 16348
rect 24232 16346 24288 16348
rect 24312 16346 24368 16348
rect 24392 16346 24448 16348
rect 24152 16294 24198 16346
rect 24198 16294 24208 16346
rect 24232 16294 24262 16346
rect 24262 16294 24274 16346
rect 24274 16294 24288 16346
rect 24312 16294 24326 16346
rect 24326 16294 24338 16346
rect 24338 16294 24368 16346
rect 24392 16294 24402 16346
rect 24402 16294 24448 16346
rect 24152 16292 24208 16294
rect 24232 16292 24288 16294
rect 24312 16292 24368 16294
rect 24392 16292 24448 16294
rect 24152 15258 24208 15260
rect 24232 15258 24288 15260
rect 24312 15258 24368 15260
rect 24392 15258 24448 15260
rect 24152 15206 24198 15258
rect 24198 15206 24208 15258
rect 24232 15206 24262 15258
rect 24262 15206 24274 15258
rect 24274 15206 24288 15258
rect 24312 15206 24326 15258
rect 24326 15206 24338 15258
rect 24338 15206 24368 15258
rect 24392 15206 24402 15258
rect 24402 15206 24448 15258
rect 24152 15204 24208 15206
rect 24232 15204 24288 15206
rect 24312 15204 24368 15206
rect 24392 15204 24448 15206
rect 23492 14714 23548 14716
rect 23572 14714 23628 14716
rect 23652 14714 23708 14716
rect 23732 14714 23788 14716
rect 23492 14662 23538 14714
rect 23538 14662 23548 14714
rect 23572 14662 23602 14714
rect 23602 14662 23614 14714
rect 23614 14662 23628 14714
rect 23652 14662 23666 14714
rect 23666 14662 23678 14714
rect 23678 14662 23708 14714
rect 23732 14662 23742 14714
rect 23742 14662 23788 14714
rect 23492 14660 23548 14662
rect 23572 14660 23628 14662
rect 23652 14660 23708 14662
rect 23732 14660 23788 14662
rect 17053 10362 17109 10364
rect 17133 10362 17189 10364
rect 17213 10362 17269 10364
rect 17293 10362 17349 10364
rect 17053 10310 17099 10362
rect 17099 10310 17109 10362
rect 17133 10310 17163 10362
rect 17163 10310 17175 10362
rect 17175 10310 17189 10362
rect 17213 10310 17227 10362
rect 17227 10310 17239 10362
rect 17239 10310 17269 10362
rect 17293 10310 17303 10362
rect 17303 10310 17349 10362
rect 17053 10308 17109 10310
rect 17133 10308 17189 10310
rect 17213 10308 17269 10310
rect 17293 10308 17349 10310
rect 17713 9818 17769 9820
rect 17793 9818 17849 9820
rect 17873 9818 17929 9820
rect 17953 9818 18009 9820
rect 17713 9766 17759 9818
rect 17759 9766 17769 9818
rect 17793 9766 17823 9818
rect 17823 9766 17835 9818
rect 17835 9766 17849 9818
rect 17873 9766 17887 9818
rect 17887 9766 17899 9818
rect 17899 9766 17929 9818
rect 17953 9766 17963 9818
rect 17963 9766 18009 9818
rect 17713 9764 17769 9766
rect 17793 9764 17849 9766
rect 17873 9764 17929 9766
rect 17953 9764 18009 9766
rect 23492 13626 23548 13628
rect 23572 13626 23628 13628
rect 23652 13626 23708 13628
rect 23732 13626 23788 13628
rect 23492 13574 23538 13626
rect 23538 13574 23548 13626
rect 23572 13574 23602 13626
rect 23602 13574 23614 13626
rect 23614 13574 23628 13626
rect 23652 13574 23666 13626
rect 23666 13574 23678 13626
rect 23678 13574 23708 13626
rect 23732 13574 23742 13626
rect 23742 13574 23788 13626
rect 23492 13572 23548 13574
rect 23572 13572 23628 13574
rect 23652 13572 23708 13574
rect 23732 13572 23788 13574
rect 24152 14170 24208 14172
rect 24232 14170 24288 14172
rect 24312 14170 24368 14172
rect 24392 14170 24448 14172
rect 24152 14118 24198 14170
rect 24198 14118 24208 14170
rect 24232 14118 24262 14170
rect 24262 14118 24274 14170
rect 24274 14118 24288 14170
rect 24312 14118 24326 14170
rect 24326 14118 24338 14170
rect 24338 14118 24368 14170
rect 24392 14118 24402 14170
rect 24402 14118 24448 14170
rect 24152 14116 24208 14118
rect 24232 14116 24288 14118
rect 24312 14116 24368 14118
rect 24392 14116 24448 14118
rect 24152 13082 24208 13084
rect 24232 13082 24288 13084
rect 24312 13082 24368 13084
rect 24392 13082 24448 13084
rect 24152 13030 24198 13082
rect 24198 13030 24208 13082
rect 24232 13030 24262 13082
rect 24262 13030 24274 13082
rect 24274 13030 24288 13082
rect 24312 13030 24326 13082
rect 24326 13030 24338 13082
rect 24338 13030 24368 13082
rect 24392 13030 24402 13082
rect 24402 13030 24448 13082
rect 24152 13028 24208 13030
rect 24232 13028 24288 13030
rect 24312 13028 24368 13030
rect 24392 13028 24448 13030
rect 23492 12538 23548 12540
rect 23572 12538 23628 12540
rect 23652 12538 23708 12540
rect 23732 12538 23788 12540
rect 23492 12486 23538 12538
rect 23538 12486 23548 12538
rect 23572 12486 23602 12538
rect 23602 12486 23614 12538
rect 23614 12486 23628 12538
rect 23652 12486 23666 12538
rect 23666 12486 23678 12538
rect 23678 12486 23708 12538
rect 23732 12486 23742 12538
rect 23742 12486 23788 12538
rect 23492 12484 23548 12486
rect 23572 12484 23628 12486
rect 23652 12484 23708 12486
rect 23732 12484 23788 12486
rect 24152 11994 24208 11996
rect 24232 11994 24288 11996
rect 24312 11994 24368 11996
rect 24392 11994 24448 11996
rect 24152 11942 24198 11994
rect 24198 11942 24208 11994
rect 24232 11942 24262 11994
rect 24262 11942 24274 11994
rect 24274 11942 24288 11994
rect 24312 11942 24326 11994
rect 24326 11942 24338 11994
rect 24338 11942 24368 11994
rect 24392 11942 24402 11994
rect 24402 11942 24448 11994
rect 24152 11940 24208 11942
rect 24232 11940 24288 11942
rect 24312 11940 24368 11942
rect 24392 11940 24448 11942
rect 23492 11450 23548 11452
rect 23572 11450 23628 11452
rect 23652 11450 23708 11452
rect 23732 11450 23788 11452
rect 23492 11398 23538 11450
rect 23538 11398 23548 11450
rect 23572 11398 23602 11450
rect 23602 11398 23614 11450
rect 23614 11398 23628 11450
rect 23652 11398 23666 11450
rect 23666 11398 23678 11450
rect 23678 11398 23708 11450
rect 23732 11398 23742 11450
rect 23742 11398 23788 11450
rect 23492 11396 23548 11398
rect 23572 11396 23628 11398
rect 23652 11396 23708 11398
rect 23732 11396 23788 11398
rect 24152 10906 24208 10908
rect 24232 10906 24288 10908
rect 24312 10906 24368 10908
rect 24392 10906 24448 10908
rect 24152 10854 24198 10906
rect 24198 10854 24208 10906
rect 24232 10854 24262 10906
rect 24262 10854 24274 10906
rect 24274 10854 24288 10906
rect 24312 10854 24326 10906
rect 24326 10854 24338 10906
rect 24338 10854 24368 10906
rect 24392 10854 24402 10906
rect 24402 10854 24448 10906
rect 24152 10852 24208 10854
rect 24232 10852 24288 10854
rect 24312 10852 24368 10854
rect 24392 10852 24448 10854
rect 23492 10362 23548 10364
rect 23572 10362 23628 10364
rect 23652 10362 23708 10364
rect 23732 10362 23788 10364
rect 23492 10310 23538 10362
rect 23538 10310 23548 10362
rect 23572 10310 23602 10362
rect 23602 10310 23614 10362
rect 23614 10310 23628 10362
rect 23652 10310 23666 10362
rect 23666 10310 23678 10362
rect 23678 10310 23708 10362
rect 23732 10310 23742 10362
rect 23742 10310 23788 10362
rect 23492 10308 23548 10310
rect 23572 10308 23628 10310
rect 23652 10308 23708 10310
rect 23732 10308 23788 10310
rect 24152 9818 24208 9820
rect 24232 9818 24288 9820
rect 24312 9818 24368 9820
rect 24392 9818 24448 9820
rect 24152 9766 24198 9818
rect 24198 9766 24208 9818
rect 24232 9766 24262 9818
rect 24262 9766 24274 9818
rect 24274 9766 24288 9818
rect 24312 9766 24326 9818
rect 24326 9766 24338 9818
rect 24338 9766 24368 9818
rect 24392 9766 24402 9818
rect 24402 9766 24448 9818
rect 24152 9764 24208 9766
rect 24232 9764 24288 9766
rect 24312 9764 24368 9766
rect 24392 9764 24448 9766
rect 17053 9274 17109 9276
rect 17133 9274 17189 9276
rect 17213 9274 17269 9276
rect 17293 9274 17349 9276
rect 17053 9222 17099 9274
rect 17099 9222 17109 9274
rect 17133 9222 17163 9274
rect 17163 9222 17175 9274
rect 17175 9222 17189 9274
rect 17213 9222 17227 9274
rect 17227 9222 17239 9274
rect 17239 9222 17269 9274
rect 17293 9222 17303 9274
rect 17303 9222 17349 9274
rect 17053 9220 17109 9222
rect 17133 9220 17189 9222
rect 17213 9220 17269 9222
rect 17293 9220 17349 9222
rect 17713 8730 17769 8732
rect 17793 8730 17849 8732
rect 17873 8730 17929 8732
rect 17953 8730 18009 8732
rect 17713 8678 17759 8730
rect 17759 8678 17769 8730
rect 17793 8678 17823 8730
rect 17823 8678 17835 8730
rect 17835 8678 17849 8730
rect 17873 8678 17887 8730
rect 17887 8678 17899 8730
rect 17899 8678 17929 8730
rect 17953 8678 17963 8730
rect 17963 8678 18009 8730
rect 17713 8676 17769 8678
rect 17793 8676 17849 8678
rect 17873 8676 17929 8678
rect 17953 8676 18009 8678
rect 17053 8186 17109 8188
rect 17133 8186 17189 8188
rect 17213 8186 17269 8188
rect 17293 8186 17349 8188
rect 17053 8134 17099 8186
rect 17099 8134 17109 8186
rect 17133 8134 17163 8186
rect 17163 8134 17175 8186
rect 17175 8134 17189 8186
rect 17213 8134 17227 8186
rect 17227 8134 17239 8186
rect 17239 8134 17269 8186
rect 17293 8134 17303 8186
rect 17303 8134 17349 8186
rect 17053 8132 17109 8134
rect 17133 8132 17189 8134
rect 17213 8132 17269 8134
rect 17293 8132 17349 8134
rect 17038 7248 17094 7304
rect 17053 7098 17109 7100
rect 17133 7098 17189 7100
rect 17213 7098 17269 7100
rect 17293 7098 17349 7100
rect 17053 7046 17099 7098
rect 17099 7046 17109 7098
rect 17133 7046 17163 7098
rect 17163 7046 17175 7098
rect 17175 7046 17189 7098
rect 17213 7046 17227 7098
rect 17227 7046 17239 7098
rect 17239 7046 17269 7098
rect 17293 7046 17303 7098
rect 17303 7046 17349 7098
rect 17053 7044 17109 7046
rect 17133 7044 17189 7046
rect 17213 7044 17269 7046
rect 17293 7044 17349 7046
rect 17713 7642 17769 7644
rect 17793 7642 17849 7644
rect 17873 7642 17929 7644
rect 17953 7642 18009 7644
rect 17713 7590 17759 7642
rect 17759 7590 17769 7642
rect 17793 7590 17823 7642
rect 17823 7590 17835 7642
rect 17835 7590 17849 7642
rect 17873 7590 17887 7642
rect 17887 7590 17899 7642
rect 17899 7590 17929 7642
rect 17953 7590 17963 7642
rect 17963 7590 18009 7642
rect 17713 7588 17769 7590
rect 17793 7588 17849 7590
rect 17873 7588 17929 7590
rect 17953 7588 18009 7590
rect 17713 6554 17769 6556
rect 17793 6554 17849 6556
rect 17873 6554 17929 6556
rect 17953 6554 18009 6556
rect 17713 6502 17759 6554
rect 17759 6502 17769 6554
rect 17793 6502 17823 6554
rect 17823 6502 17835 6554
rect 17835 6502 17849 6554
rect 17873 6502 17887 6554
rect 17887 6502 17899 6554
rect 17899 6502 17929 6554
rect 17953 6502 17963 6554
rect 17963 6502 18009 6554
rect 17713 6500 17769 6502
rect 17793 6500 17849 6502
rect 17873 6500 17929 6502
rect 17953 6500 18009 6502
rect 17053 6010 17109 6012
rect 17133 6010 17189 6012
rect 17213 6010 17269 6012
rect 17293 6010 17349 6012
rect 17053 5958 17099 6010
rect 17099 5958 17109 6010
rect 17133 5958 17163 6010
rect 17163 5958 17175 6010
rect 17175 5958 17189 6010
rect 17213 5958 17227 6010
rect 17227 5958 17239 6010
rect 17239 5958 17269 6010
rect 17293 5958 17303 6010
rect 17303 5958 17349 6010
rect 17053 5956 17109 5958
rect 17133 5956 17189 5958
rect 17213 5956 17269 5958
rect 17293 5956 17349 5958
rect 17713 5466 17769 5468
rect 17793 5466 17849 5468
rect 17873 5466 17929 5468
rect 17953 5466 18009 5468
rect 17713 5414 17759 5466
rect 17759 5414 17769 5466
rect 17793 5414 17823 5466
rect 17823 5414 17835 5466
rect 17835 5414 17849 5466
rect 17873 5414 17887 5466
rect 17887 5414 17899 5466
rect 17899 5414 17929 5466
rect 17953 5414 17963 5466
rect 17963 5414 18009 5466
rect 17713 5412 17769 5414
rect 17793 5412 17849 5414
rect 17873 5412 17929 5414
rect 17953 5412 18009 5414
rect 17053 4922 17109 4924
rect 17133 4922 17189 4924
rect 17213 4922 17269 4924
rect 17293 4922 17349 4924
rect 17053 4870 17099 4922
rect 17099 4870 17109 4922
rect 17133 4870 17163 4922
rect 17163 4870 17175 4922
rect 17175 4870 17189 4922
rect 17213 4870 17227 4922
rect 17227 4870 17239 4922
rect 17239 4870 17269 4922
rect 17293 4870 17303 4922
rect 17303 4870 17349 4922
rect 17053 4868 17109 4870
rect 17133 4868 17189 4870
rect 17213 4868 17269 4870
rect 17293 4868 17349 4870
rect 16762 4392 16818 4448
rect 17713 4378 17769 4380
rect 17793 4378 17849 4380
rect 17873 4378 17929 4380
rect 17953 4378 18009 4380
rect 17713 4326 17759 4378
rect 17759 4326 17769 4378
rect 17793 4326 17823 4378
rect 17823 4326 17835 4378
rect 17835 4326 17849 4378
rect 17873 4326 17887 4378
rect 17887 4326 17899 4378
rect 17899 4326 17929 4378
rect 17953 4326 17963 4378
rect 17963 4326 18009 4378
rect 17713 4324 17769 4326
rect 17793 4324 17849 4326
rect 17873 4324 17929 4326
rect 17953 4324 18009 4326
rect 17774 3984 17830 4040
rect 17053 3834 17109 3836
rect 17133 3834 17189 3836
rect 17213 3834 17269 3836
rect 17293 3834 17349 3836
rect 17053 3782 17099 3834
rect 17099 3782 17109 3834
rect 17133 3782 17163 3834
rect 17163 3782 17175 3834
rect 17175 3782 17189 3834
rect 17213 3782 17227 3834
rect 17227 3782 17239 3834
rect 17239 3782 17269 3834
rect 17293 3782 17303 3834
rect 17303 3782 17349 3834
rect 17053 3780 17109 3782
rect 17133 3780 17189 3782
rect 17213 3780 17269 3782
rect 17293 3780 17349 3782
rect 23492 9274 23548 9276
rect 23572 9274 23628 9276
rect 23652 9274 23708 9276
rect 23732 9274 23788 9276
rect 23492 9222 23538 9274
rect 23538 9222 23548 9274
rect 23572 9222 23602 9274
rect 23602 9222 23614 9274
rect 23614 9222 23628 9274
rect 23652 9222 23666 9274
rect 23666 9222 23678 9274
rect 23678 9222 23708 9274
rect 23732 9222 23742 9274
rect 23742 9222 23788 9274
rect 23492 9220 23548 9222
rect 23572 9220 23628 9222
rect 23652 9220 23708 9222
rect 23732 9220 23788 9222
rect 24152 8730 24208 8732
rect 24232 8730 24288 8732
rect 24312 8730 24368 8732
rect 24392 8730 24448 8732
rect 24152 8678 24198 8730
rect 24198 8678 24208 8730
rect 24232 8678 24262 8730
rect 24262 8678 24274 8730
rect 24274 8678 24288 8730
rect 24312 8678 24326 8730
rect 24326 8678 24338 8730
rect 24338 8678 24368 8730
rect 24392 8678 24402 8730
rect 24402 8678 24448 8730
rect 24152 8676 24208 8678
rect 24232 8676 24288 8678
rect 24312 8676 24368 8678
rect 24392 8676 24448 8678
rect 26514 11192 26570 11248
rect 23492 8186 23548 8188
rect 23572 8186 23628 8188
rect 23652 8186 23708 8188
rect 23732 8186 23788 8188
rect 23492 8134 23538 8186
rect 23538 8134 23548 8186
rect 23572 8134 23602 8186
rect 23602 8134 23614 8186
rect 23614 8134 23628 8186
rect 23652 8134 23666 8186
rect 23666 8134 23678 8186
rect 23678 8134 23708 8186
rect 23732 8134 23742 8186
rect 23742 8134 23788 8186
rect 23492 8132 23548 8134
rect 23572 8132 23628 8134
rect 23652 8132 23708 8134
rect 23732 8132 23788 8134
rect 24152 7642 24208 7644
rect 24232 7642 24288 7644
rect 24312 7642 24368 7644
rect 24392 7642 24448 7644
rect 24152 7590 24198 7642
rect 24198 7590 24208 7642
rect 24232 7590 24262 7642
rect 24262 7590 24274 7642
rect 24274 7590 24288 7642
rect 24312 7590 24326 7642
rect 24326 7590 24338 7642
rect 24338 7590 24368 7642
rect 24392 7590 24402 7642
rect 24402 7590 24448 7642
rect 24152 7588 24208 7590
rect 24232 7588 24288 7590
rect 24312 7588 24368 7590
rect 24392 7588 24448 7590
rect 25686 7384 25742 7440
rect 23492 7098 23548 7100
rect 23572 7098 23628 7100
rect 23652 7098 23708 7100
rect 23732 7098 23788 7100
rect 23492 7046 23538 7098
rect 23538 7046 23548 7098
rect 23572 7046 23602 7098
rect 23602 7046 23614 7098
rect 23614 7046 23628 7098
rect 23652 7046 23666 7098
rect 23666 7046 23678 7098
rect 23678 7046 23708 7098
rect 23732 7046 23742 7098
rect 23742 7046 23788 7098
rect 23492 7044 23548 7046
rect 23572 7044 23628 7046
rect 23652 7044 23708 7046
rect 23732 7044 23788 7046
rect 24152 6554 24208 6556
rect 24232 6554 24288 6556
rect 24312 6554 24368 6556
rect 24392 6554 24448 6556
rect 24152 6502 24198 6554
rect 24198 6502 24208 6554
rect 24232 6502 24262 6554
rect 24262 6502 24274 6554
rect 24274 6502 24288 6554
rect 24312 6502 24326 6554
rect 24326 6502 24338 6554
rect 24338 6502 24368 6554
rect 24392 6502 24402 6554
rect 24402 6502 24448 6554
rect 24152 6500 24208 6502
rect 24232 6500 24288 6502
rect 24312 6500 24368 6502
rect 24392 6500 24448 6502
rect 23492 6010 23548 6012
rect 23572 6010 23628 6012
rect 23652 6010 23708 6012
rect 23732 6010 23788 6012
rect 23492 5958 23538 6010
rect 23538 5958 23548 6010
rect 23572 5958 23602 6010
rect 23602 5958 23614 6010
rect 23614 5958 23628 6010
rect 23652 5958 23666 6010
rect 23666 5958 23678 6010
rect 23678 5958 23708 6010
rect 23732 5958 23742 6010
rect 23742 5958 23788 6010
rect 23492 5956 23548 5958
rect 23572 5956 23628 5958
rect 23652 5956 23708 5958
rect 23732 5956 23788 5958
rect 24152 5466 24208 5468
rect 24232 5466 24288 5468
rect 24312 5466 24368 5468
rect 24392 5466 24448 5468
rect 24152 5414 24198 5466
rect 24198 5414 24208 5466
rect 24232 5414 24262 5466
rect 24262 5414 24274 5466
rect 24274 5414 24288 5466
rect 24312 5414 24326 5466
rect 24326 5414 24338 5466
rect 24338 5414 24368 5466
rect 24392 5414 24402 5466
rect 24402 5414 24448 5466
rect 24152 5412 24208 5414
rect 24232 5412 24288 5414
rect 24312 5412 24368 5414
rect 24392 5412 24448 5414
rect 23492 4922 23548 4924
rect 23572 4922 23628 4924
rect 23652 4922 23708 4924
rect 23732 4922 23788 4924
rect 23492 4870 23538 4922
rect 23538 4870 23548 4922
rect 23572 4870 23602 4922
rect 23602 4870 23614 4922
rect 23614 4870 23628 4922
rect 23652 4870 23666 4922
rect 23666 4870 23678 4922
rect 23678 4870 23708 4922
rect 23732 4870 23742 4922
rect 23742 4870 23788 4922
rect 23492 4868 23548 4870
rect 23572 4868 23628 4870
rect 23652 4868 23708 4870
rect 23732 4868 23788 4870
rect 24152 4378 24208 4380
rect 24232 4378 24288 4380
rect 24312 4378 24368 4380
rect 24392 4378 24448 4380
rect 24152 4326 24198 4378
rect 24198 4326 24208 4378
rect 24232 4326 24262 4378
rect 24262 4326 24274 4378
rect 24274 4326 24288 4378
rect 24312 4326 24326 4378
rect 24326 4326 24338 4378
rect 24338 4326 24368 4378
rect 24392 4326 24402 4378
rect 24402 4326 24448 4378
rect 24152 4324 24208 4326
rect 24232 4324 24288 4326
rect 24312 4324 24368 4326
rect 24392 4324 24448 4326
rect 17713 3290 17769 3292
rect 17793 3290 17849 3292
rect 17873 3290 17929 3292
rect 17953 3290 18009 3292
rect 17713 3238 17759 3290
rect 17759 3238 17769 3290
rect 17793 3238 17823 3290
rect 17823 3238 17835 3290
rect 17835 3238 17849 3290
rect 17873 3238 17887 3290
rect 17887 3238 17899 3290
rect 17899 3238 17929 3290
rect 17953 3238 17963 3290
rect 17963 3238 18009 3290
rect 17713 3236 17769 3238
rect 17793 3236 17849 3238
rect 17873 3236 17929 3238
rect 17953 3236 18009 3238
rect 26514 3848 26570 3904
rect 23492 3834 23548 3836
rect 23572 3834 23628 3836
rect 23652 3834 23708 3836
rect 23732 3834 23788 3836
rect 23492 3782 23538 3834
rect 23538 3782 23548 3834
rect 23572 3782 23602 3834
rect 23602 3782 23614 3834
rect 23614 3782 23628 3834
rect 23652 3782 23666 3834
rect 23666 3782 23678 3834
rect 23678 3782 23708 3834
rect 23732 3782 23742 3834
rect 23742 3782 23788 3834
rect 23492 3780 23548 3782
rect 23572 3780 23628 3782
rect 23652 3780 23708 3782
rect 23732 3780 23788 3782
rect 24152 3290 24208 3292
rect 24232 3290 24288 3292
rect 24312 3290 24368 3292
rect 24392 3290 24448 3292
rect 24152 3238 24198 3290
rect 24198 3238 24208 3290
rect 24232 3238 24262 3290
rect 24262 3238 24274 3290
rect 24274 3238 24288 3290
rect 24312 3238 24326 3290
rect 24326 3238 24338 3290
rect 24338 3238 24368 3290
rect 24392 3238 24402 3290
rect 24402 3238 24448 3290
rect 24152 3236 24208 3238
rect 24232 3236 24288 3238
rect 24312 3236 24368 3238
rect 24392 3236 24448 3238
rect 17053 2746 17109 2748
rect 17133 2746 17189 2748
rect 17213 2746 17269 2748
rect 17293 2746 17349 2748
rect 17053 2694 17099 2746
rect 17099 2694 17109 2746
rect 17133 2694 17163 2746
rect 17163 2694 17175 2746
rect 17175 2694 17189 2746
rect 17213 2694 17227 2746
rect 17227 2694 17239 2746
rect 17239 2694 17269 2746
rect 17293 2694 17303 2746
rect 17303 2694 17349 2746
rect 17053 2692 17109 2694
rect 17133 2692 17189 2694
rect 17213 2692 17269 2694
rect 17293 2692 17349 2694
rect 23492 2746 23548 2748
rect 23572 2746 23628 2748
rect 23652 2746 23708 2748
rect 23732 2746 23788 2748
rect 23492 2694 23538 2746
rect 23538 2694 23548 2746
rect 23572 2694 23602 2746
rect 23602 2694 23614 2746
rect 23614 2694 23628 2746
rect 23652 2694 23666 2746
rect 23666 2694 23678 2746
rect 23678 2694 23708 2746
rect 23732 2694 23742 2746
rect 23742 2694 23788 2746
rect 23492 2692 23548 2694
rect 23572 2692 23628 2694
rect 23652 2692 23708 2694
rect 23732 2692 23788 2694
rect 4835 2202 4891 2204
rect 4915 2202 4971 2204
rect 4995 2202 5051 2204
rect 5075 2202 5131 2204
rect 4835 2150 4881 2202
rect 4881 2150 4891 2202
rect 4915 2150 4945 2202
rect 4945 2150 4957 2202
rect 4957 2150 4971 2202
rect 4995 2150 5009 2202
rect 5009 2150 5021 2202
rect 5021 2150 5051 2202
rect 5075 2150 5085 2202
rect 5085 2150 5131 2202
rect 4835 2148 4891 2150
rect 4915 2148 4971 2150
rect 4995 2148 5051 2150
rect 5075 2148 5131 2150
rect 11274 2202 11330 2204
rect 11354 2202 11410 2204
rect 11434 2202 11490 2204
rect 11514 2202 11570 2204
rect 11274 2150 11320 2202
rect 11320 2150 11330 2202
rect 11354 2150 11384 2202
rect 11384 2150 11396 2202
rect 11396 2150 11410 2202
rect 11434 2150 11448 2202
rect 11448 2150 11460 2202
rect 11460 2150 11490 2202
rect 11514 2150 11524 2202
rect 11524 2150 11570 2202
rect 11274 2148 11330 2150
rect 11354 2148 11410 2150
rect 11434 2148 11490 2150
rect 11514 2148 11570 2150
rect 17713 2202 17769 2204
rect 17793 2202 17849 2204
rect 17873 2202 17929 2204
rect 17953 2202 18009 2204
rect 17713 2150 17759 2202
rect 17759 2150 17769 2202
rect 17793 2150 17823 2202
rect 17823 2150 17835 2202
rect 17835 2150 17849 2202
rect 17873 2150 17887 2202
rect 17887 2150 17899 2202
rect 17899 2150 17929 2202
rect 17953 2150 17963 2202
rect 17963 2150 18009 2202
rect 17713 2148 17769 2150
rect 17793 2148 17849 2150
rect 17873 2148 17929 2150
rect 17953 2148 18009 2150
rect 24152 2202 24208 2204
rect 24232 2202 24288 2204
rect 24312 2202 24368 2204
rect 24392 2202 24448 2204
rect 24152 2150 24198 2202
rect 24198 2150 24208 2202
rect 24232 2150 24262 2202
rect 24262 2150 24274 2202
rect 24274 2150 24288 2202
rect 24312 2150 24326 2202
rect 24326 2150 24338 2202
rect 24338 2150 24368 2202
rect 24392 2150 24402 2202
rect 24402 2150 24448 2202
rect 24152 2148 24208 2150
rect 24232 2148 24288 2150
rect 24312 2148 24368 2150
rect 24392 2148 24448 2150
<< metal3 >>
rect 0 28114 800 28144
rect 2221 28114 2287 28117
rect 0 28112 2287 28114
rect 0 28056 2226 28112
rect 2282 28056 2287 28112
rect 0 28054 2287 28056
rect 0 28024 800 28054
rect 2221 28051 2287 28054
rect 4165 27776 4481 27777
rect 4165 27712 4171 27776
rect 4235 27712 4251 27776
rect 4315 27712 4331 27776
rect 4395 27712 4411 27776
rect 4475 27712 4481 27776
rect 4165 27711 4481 27712
rect 10604 27776 10920 27777
rect 10604 27712 10610 27776
rect 10674 27712 10690 27776
rect 10754 27712 10770 27776
rect 10834 27712 10850 27776
rect 10914 27712 10920 27776
rect 10604 27711 10920 27712
rect 17043 27776 17359 27777
rect 17043 27712 17049 27776
rect 17113 27712 17129 27776
rect 17193 27712 17209 27776
rect 17273 27712 17289 27776
rect 17353 27712 17359 27776
rect 17043 27711 17359 27712
rect 23482 27776 23798 27777
rect 23482 27712 23488 27776
rect 23552 27712 23568 27776
rect 23632 27712 23648 27776
rect 23712 27712 23728 27776
rect 23792 27712 23798 27776
rect 23482 27711 23798 27712
rect 4825 27232 5141 27233
rect 4825 27168 4831 27232
rect 4895 27168 4911 27232
rect 4975 27168 4991 27232
rect 5055 27168 5071 27232
rect 5135 27168 5141 27232
rect 4825 27167 5141 27168
rect 11264 27232 11580 27233
rect 11264 27168 11270 27232
rect 11334 27168 11350 27232
rect 11414 27168 11430 27232
rect 11494 27168 11510 27232
rect 11574 27168 11580 27232
rect 11264 27167 11580 27168
rect 17703 27232 18019 27233
rect 17703 27168 17709 27232
rect 17773 27168 17789 27232
rect 17853 27168 17869 27232
rect 17933 27168 17949 27232
rect 18013 27168 18019 27232
rect 17703 27167 18019 27168
rect 24142 27232 24458 27233
rect 24142 27168 24148 27232
rect 24212 27168 24228 27232
rect 24292 27168 24308 27232
rect 24372 27168 24388 27232
rect 24452 27168 24458 27232
rect 24142 27167 24458 27168
rect 4165 26688 4481 26689
rect 4165 26624 4171 26688
rect 4235 26624 4251 26688
rect 4315 26624 4331 26688
rect 4395 26624 4411 26688
rect 4475 26624 4481 26688
rect 4165 26623 4481 26624
rect 10604 26688 10920 26689
rect 10604 26624 10610 26688
rect 10674 26624 10690 26688
rect 10754 26624 10770 26688
rect 10834 26624 10850 26688
rect 10914 26624 10920 26688
rect 10604 26623 10920 26624
rect 17043 26688 17359 26689
rect 17043 26624 17049 26688
rect 17113 26624 17129 26688
rect 17193 26624 17209 26688
rect 17273 26624 17289 26688
rect 17353 26624 17359 26688
rect 17043 26623 17359 26624
rect 23482 26688 23798 26689
rect 23482 26624 23488 26688
rect 23552 26624 23568 26688
rect 23632 26624 23648 26688
rect 23712 26624 23728 26688
rect 23792 26624 23798 26688
rect 23482 26623 23798 26624
rect 4825 26144 5141 26145
rect 4825 26080 4831 26144
rect 4895 26080 4911 26144
rect 4975 26080 4991 26144
rect 5055 26080 5071 26144
rect 5135 26080 5141 26144
rect 4825 26079 5141 26080
rect 11264 26144 11580 26145
rect 11264 26080 11270 26144
rect 11334 26080 11350 26144
rect 11414 26080 11430 26144
rect 11494 26080 11510 26144
rect 11574 26080 11580 26144
rect 11264 26079 11580 26080
rect 17703 26144 18019 26145
rect 17703 26080 17709 26144
rect 17773 26080 17789 26144
rect 17853 26080 17869 26144
rect 17933 26080 17949 26144
rect 18013 26080 18019 26144
rect 17703 26079 18019 26080
rect 24142 26144 24458 26145
rect 24142 26080 24148 26144
rect 24212 26080 24228 26144
rect 24292 26080 24308 26144
rect 24372 26080 24388 26144
rect 24452 26080 24458 26144
rect 24142 26079 24458 26080
rect 0 25938 800 25968
rect 3417 25938 3483 25941
rect 0 25936 3483 25938
rect 0 25880 3422 25936
rect 3478 25880 3483 25936
rect 0 25878 3483 25880
rect 0 25848 800 25878
rect 3417 25875 3483 25878
rect 26141 25938 26207 25941
rect 27188 25938 27988 25968
rect 26141 25936 27988 25938
rect 26141 25880 26146 25936
rect 26202 25880 27988 25936
rect 26141 25878 27988 25880
rect 26141 25875 26207 25878
rect 27188 25848 27988 25878
rect 4165 25600 4481 25601
rect 4165 25536 4171 25600
rect 4235 25536 4251 25600
rect 4315 25536 4331 25600
rect 4395 25536 4411 25600
rect 4475 25536 4481 25600
rect 4165 25535 4481 25536
rect 10604 25600 10920 25601
rect 10604 25536 10610 25600
rect 10674 25536 10690 25600
rect 10754 25536 10770 25600
rect 10834 25536 10850 25600
rect 10914 25536 10920 25600
rect 10604 25535 10920 25536
rect 17043 25600 17359 25601
rect 17043 25536 17049 25600
rect 17113 25536 17129 25600
rect 17193 25536 17209 25600
rect 17273 25536 17289 25600
rect 17353 25536 17359 25600
rect 17043 25535 17359 25536
rect 23482 25600 23798 25601
rect 23482 25536 23488 25600
rect 23552 25536 23568 25600
rect 23632 25536 23648 25600
rect 23712 25536 23728 25600
rect 23792 25536 23798 25600
rect 23482 25535 23798 25536
rect 4825 25056 5141 25057
rect 4825 24992 4831 25056
rect 4895 24992 4911 25056
rect 4975 24992 4991 25056
rect 5055 24992 5071 25056
rect 5135 24992 5141 25056
rect 4825 24991 5141 24992
rect 11264 25056 11580 25057
rect 11264 24992 11270 25056
rect 11334 24992 11350 25056
rect 11414 24992 11430 25056
rect 11494 24992 11510 25056
rect 11574 24992 11580 25056
rect 11264 24991 11580 24992
rect 17703 25056 18019 25057
rect 17703 24992 17709 25056
rect 17773 24992 17789 25056
rect 17853 24992 17869 25056
rect 17933 24992 17949 25056
rect 18013 24992 18019 25056
rect 17703 24991 18019 24992
rect 24142 25056 24458 25057
rect 24142 24992 24148 25056
rect 24212 24992 24228 25056
rect 24292 24992 24308 25056
rect 24372 24992 24388 25056
rect 24452 24992 24458 25056
rect 24142 24991 24458 24992
rect 4165 24512 4481 24513
rect 4165 24448 4171 24512
rect 4235 24448 4251 24512
rect 4315 24448 4331 24512
rect 4395 24448 4411 24512
rect 4475 24448 4481 24512
rect 4165 24447 4481 24448
rect 10604 24512 10920 24513
rect 10604 24448 10610 24512
rect 10674 24448 10690 24512
rect 10754 24448 10770 24512
rect 10834 24448 10850 24512
rect 10914 24448 10920 24512
rect 10604 24447 10920 24448
rect 17043 24512 17359 24513
rect 17043 24448 17049 24512
rect 17113 24448 17129 24512
rect 17193 24448 17209 24512
rect 17273 24448 17289 24512
rect 17353 24448 17359 24512
rect 17043 24447 17359 24448
rect 23482 24512 23798 24513
rect 23482 24448 23488 24512
rect 23552 24448 23568 24512
rect 23632 24448 23648 24512
rect 23712 24448 23728 24512
rect 23792 24448 23798 24512
rect 23482 24447 23798 24448
rect 4825 23968 5141 23969
rect 4825 23904 4831 23968
rect 4895 23904 4911 23968
rect 4975 23904 4991 23968
rect 5055 23904 5071 23968
rect 5135 23904 5141 23968
rect 4825 23903 5141 23904
rect 11264 23968 11580 23969
rect 11264 23904 11270 23968
rect 11334 23904 11350 23968
rect 11414 23904 11430 23968
rect 11494 23904 11510 23968
rect 11574 23904 11580 23968
rect 11264 23903 11580 23904
rect 17703 23968 18019 23969
rect 17703 23904 17709 23968
rect 17773 23904 17789 23968
rect 17853 23904 17869 23968
rect 17933 23904 17949 23968
rect 18013 23904 18019 23968
rect 17703 23903 18019 23904
rect 24142 23968 24458 23969
rect 24142 23904 24148 23968
rect 24212 23904 24228 23968
rect 24292 23904 24308 23968
rect 24372 23904 24388 23968
rect 24452 23904 24458 23968
rect 24142 23903 24458 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 9305 23762 9371 23765
rect 10317 23762 10383 23765
rect 9305 23760 10383 23762
rect 9305 23704 9310 23760
rect 9366 23704 10322 23760
rect 10378 23704 10383 23760
rect 9305 23702 10383 23704
rect 9305 23699 9371 23702
rect 10317 23699 10383 23702
rect 9765 23626 9831 23629
rect 10593 23626 10659 23629
rect 9765 23624 10659 23626
rect 9765 23568 9770 23624
rect 9826 23568 10598 23624
rect 10654 23568 10659 23624
rect 9765 23566 10659 23568
rect 9765 23563 9831 23566
rect 10593 23563 10659 23566
rect 4165 23424 4481 23425
rect 4165 23360 4171 23424
rect 4235 23360 4251 23424
rect 4315 23360 4331 23424
rect 4395 23360 4411 23424
rect 4475 23360 4481 23424
rect 4165 23359 4481 23360
rect 10604 23424 10920 23425
rect 10604 23360 10610 23424
rect 10674 23360 10690 23424
rect 10754 23360 10770 23424
rect 10834 23360 10850 23424
rect 10914 23360 10920 23424
rect 10604 23359 10920 23360
rect 17043 23424 17359 23425
rect 17043 23360 17049 23424
rect 17113 23360 17129 23424
rect 17193 23360 17209 23424
rect 17273 23360 17289 23424
rect 17353 23360 17359 23424
rect 17043 23359 17359 23360
rect 23482 23424 23798 23425
rect 23482 23360 23488 23424
rect 23552 23360 23568 23424
rect 23632 23360 23648 23424
rect 23712 23360 23728 23424
rect 23792 23360 23798 23424
rect 23482 23359 23798 23360
rect 9029 23354 9095 23357
rect 9857 23354 9923 23357
rect 9029 23352 9923 23354
rect 9029 23296 9034 23352
rect 9090 23296 9862 23352
rect 9918 23296 9923 23352
rect 9029 23294 9923 23296
rect 9029 23291 9095 23294
rect 9857 23291 9923 23294
rect 6177 23218 6243 23221
rect 15837 23218 15903 23221
rect 6177 23216 15903 23218
rect 6177 23160 6182 23216
rect 6238 23160 15842 23216
rect 15898 23160 15903 23216
rect 6177 23158 15903 23160
rect 6177 23155 6243 23158
rect 15837 23155 15903 23158
rect 8937 23082 9003 23085
rect 9765 23082 9831 23085
rect 8937 23080 9831 23082
rect 8937 23024 8942 23080
rect 8998 23024 9770 23080
rect 9826 23024 9831 23080
rect 8937 23022 9831 23024
rect 8937 23019 9003 23022
rect 9765 23019 9831 23022
rect 11421 23082 11487 23085
rect 18229 23082 18295 23085
rect 11421 23080 18295 23082
rect 11421 23024 11426 23080
rect 11482 23024 18234 23080
rect 18290 23024 18295 23080
rect 11421 23022 18295 23024
rect 11421 23019 11487 23022
rect 18229 23019 18295 23022
rect 4825 22880 5141 22881
rect 4825 22816 4831 22880
rect 4895 22816 4911 22880
rect 4975 22816 4991 22880
rect 5055 22816 5071 22880
rect 5135 22816 5141 22880
rect 4825 22815 5141 22816
rect 11264 22880 11580 22881
rect 11264 22816 11270 22880
rect 11334 22816 11350 22880
rect 11414 22816 11430 22880
rect 11494 22816 11510 22880
rect 11574 22816 11580 22880
rect 11264 22815 11580 22816
rect 17703 22880 18019 22881
rect 17703 22816 17709 22880
rect 17773 22816 17789 22880
rect 17853 22816 17869 22880
rect 17933 22816 17949 22880
rect 18013 22816 18019 22880
rect 17703 22815 18019 22816
rect 24142 22880 24458 22881
rect 24142 22816 24148 22880
rect 24212 22816 24228 22880
rect 24292 22816 24308 22880
rect 24372 22816 24388 22880
rect 24452 22816 24458 22880
rect 24142 22815 24458 22816
rect 9121 22674 9187 22677
rect 11973 22674 12039 22677
rect 9121 22672 12039 22674
rect 9121 22616 9126 22672
rect 9182 22616 11978 22672
rect 12034 22616 12039 22672
rect 9121 22614 12039 22616
rect 9121 22611 9187 22614
rect 11973 22611 12039 22614
rect 9673 22538 9739 22541
rect 12709 22538 12775 22541
rect 9673 22536 12775 22538
rect 9673 22480 9678 22536
rect 9734 22480 12714 22536
rect 12770 22480 12775 22536
rect 9673 22478 12775 22480
rect 9673 22475 9739 22478
rect 12709 22475 12775 22478
rect 4165 22336 4481 22337
rect 4165 22272 4171 22336
rect 4235 22272 4251 22336
rect 4315 22272 4331 22336
rect 4395 22272 4411 22336
rect 4475 22272 4481 22336
rect 4165 22271 4481 22272
rect 10604 22336 10920 22337
rect 10604 22272 10610 22336
rect 10674 22272 10690 22336
rect 10754 22272 10770 22336
rect 10834 22272 10850 22336
rect 10914 22272 10920 22336
rect 10604 22271 10920 22272
rect 17043 22336 17359 22337
rect 17043 22272 17049 22336
rect 17113 22272 17129 22336
rect 17193 22272 17209 22336
rect 17273 22272 17289 22336
rect 17353 22272 17359 22336
rect 17043 22271 17359 22272
rect 23482 22336 23798 22337
rect 23482 22272 23488 22336
rect 23552 22272 23568 22336
rect 23632 22272 23648 22336
rect 23712 22272 23728 22336
rect 23792 22272 23798 22336
rect 23482 22271 23798 22272
rect 11053 22130 11119 22133
rect 18045 22130 18111 22133
rect 11053 22128 18111 22130
rect 11053 22072 11058 22128
rect 11114 22072 18050 22128
rect 18106 22072 18111 22128
rect 11053 22070 18111 22072
rect 11053 22067 11119 22070
rect 18045 22067 18111 22070
rect 4061 21994 4127 21997
rect 5073 21994 5139 21997
rect 4061 21992 5139 21994
rect 4061 21936 4066 21992
rect 4122 21936 5078 21992
rect 5134 21936 5139 21992
rect 4061 21934 5139 21936
rect 4061 21931 4127 21934
rect 5073 21931 5139 21934
rect 9857 21994 9923 21997
rect 11605 21994 11671 21997
rect 9857 21992 11671 21994
rect 9857 21936 9862 21992
rect 9918 21936 11610 21992
rect 11666 21936 11671 21992
rect 9857 21934 11671 21936
rect 9857 21931 9923 21934
rect 11605 21931 11671 21934
rect 4825 21792 5141 21793
rect 4825 21728 4831 21792
rect 4895 21728 4911 21792
rect 4975 21728 4991 21792
rect 5055 21728 5071 21792
rect 5135 21728 5141 21792
rect 4825 21727 5141 21728
rect 11264 21792 11580 21793
rect 11264 21728 11270 21792
rect 11334 21728 11350 21792
rect 11414 21728 11430 21792
rect 11494 21728 11510 21792
rect 11574 21728 11580 21792
rect 11264 21727 11580 21728
rect 17703 21792 18019 21793
rect 17703 21728 17709 21792
rect 17773 21728 17789 21792
rect 17853 21728 17869 21792
rect 17933 21728 17949 21792
rect 18013 21728 18019 21792
rect 17703 21727 18019 21728
rect 24142 21792 24458 21793
rect 24142 21728 24148 21792
rect 24212 21728 24228 21792
rect 24292 21728 24308 21792
rect 24372 21728 24388 21792
rect 24452 21728 24458 21792
rect 24142 21727 24458 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 4165 21248 4481 21249
rect 4165 21184 4171 21248
rect 4235 21184 4251 21248
rect 4315 21184 4331 21248
rect 4395 21184 4411 21248
rect 4475 21184 4481 21248
rect 4165 21183 4481 21184
rect 10604 21248 10920 21249
rect 10604 21184 10610 21248
rect 10674 21184 10690 21248
rect 10754 21184 10770 21248
rect 10834 21184 10850 21248
rect 10914 21184 10920 21248
rect 10604 21183 10920 21184
rect 17043 21248 17359 21249
rect 17043 21184 17049 21248
rect 17113 21184 17129 21248
rect 17193 21184 17209 21248
rect 17273 21184 17289 21248
rect 17353 21184 17359 21248
rect 17043 21183 17359 21184
rect 23482 21248 23798 21249
rect 23482 21184 23488 21248
rect 23552 21184 23568 21248
rect 23632 21184 23648 21248
rect 23712 21184 23728 21248
rect 23792 21184 23798 21248
rect 23482 21183 23798 21184
rect 14549 20770 14615 20773
rect 15326 20770 15332 20772
rect 14549 20768 15332 20770
rect 14549 20712 14554 20768
rect 14610 20712 15332 20768
rect 14549 20710 15332 20712
rect 14549 20707 14615 20710
rect 15326 20708 15332 20710
rect 15396 20708 15402 20772
rect 4825 20704 5141 20705
rect 4825 20640 4831 20704
rect 4895 20640 4911 20704
rect 4975 20640 4991 20704
rect 5055 20640 5071 20704
rect 5135 20640 5141 20704
rect 4825 20639 5141 20640
rect 11264 20704 11580 20705
rect 11264 20640 11270 20704
rect 11334 20640 11350 20704
rect 11414 20640 11430 20704
rect 11494 20640 11510 20704
rect 11574 20640 11580 20704
rect 11264 20639 11580 20640
rect 17703 20704 18019 20705
rect 17703 20640 17709 20704
rect 17773 20640 17789 20704
rect 17853 20640 17869 20704
rect 17933 20640 17949 20704
rect 18013 20640 18019 20704
rect 17703 20639 18019 20640
rect 24142 20704 24458 20705
rect 24142 20640 24148 20704
rect 24212 20640 24228 20704
rect 24292 20640 24308 20704
rect 24372 20640 24388 20704
rect 24452 20640 24458 20704
rect 24142 20639 24458 20640
rect 15510 20436 15516 20500
rect 15580 20498 15586 20500
rect 17033 20498 17099 20501
rect 15580 20496 17099 20498
rect 15580 20440 17038 20496
rect 17094 20440 17099 20496
rect 15580 20438 17099 20440
rect 15580 20436 15586 20438
rect 17033 20435 17099 20438
rect 15837 20362 15903 20365
rect 10366 20360 15903 20362
rect 10366 20304 15842 20360
rect 15898 20304 15903 20360
rect 10366 20302 15903 20304
rect 4165 20160 4481 20161
rect 4165 20096 4171 20160
rect 4235 20096 4251 20160
rect 4315 20096 4331 20160
rect 4395 20096 4411 20160
rect 4475 20096 4481 20160
rect 4165 20095 4481 20096
rect 10366 20093 10426 20302
rect 15837 20299 15903 20302
rect 16389 20362 16455 20365
rect 25497 20362 25563 20365
rect 16389 20360 25563 20362
rect 16389 20304 16394 20360
rect 16450 20304 25502 20360
rect 25558 20304 25563 20360
rect 16389 20302 25563 20304
rect 16389 20299 16455 20302
rect 25497 20299 25563 20302
rect 10604 20160 10920 20161
rect 10604 20096 10610 20160
rect 10674 20096 10690 20160
rect 10754 20096 10770 20160
rect 10834 20096 10850 20160
rect 10914 20096 10920 20160
rect 10604 20095 10920 20096
rect 17043 20160 17359 20161
rect 17043 20096 17049 20160
rect 17113 20096 17129 20160
rect 17193 20096 17209 20160
rect 17273 20096 17289 20160
rect 17353 20096 17359 20160
rect 17043 20095 17359 20096
rect 23482 20160 23798 20161
rect 23482 20096 23488 20160
rect 23552 20096 23568 20160
rect 23632 20096 23648 20160
rect 23712 20096 23728 20160
rect 23792 20096 23798 20160
rect 23482 20095 23798 20096
rect 10317 20088 10426 20093
rect 10317 20032 10322 20088
rect 10378 20032 10426 20088
rect 10317 20030 10426 20032
rect 10317 20027 10383 20030
rect 1577 19954 1643 19957
rect 12249 19954 12315 19957
rect 1577 19952 12315 19954
rect 1577 19896 1582 19952
rect 1638 19896 12254 19952
rect 12310 19896 12315 19952
rect 1577 19894 12315 19896
rect 1577 19891 1643 19894
rect 12249 19891 12315 19894
rect 1577 19818 1643 19821
rect 11789 19818 11855 19821
rect 1577 19816 11855 19818
rect 1577 19760 1582 19816
rect 1638 19760 11794 19816
rect 11850 19760 11855 19816
rect 1577 19758 11855 19760
rect 1577 19755 1643 19758
rect 11789 19755 11855 19758
rect 4825 19616 5141 19617
rect 4825 19552 4831 19616
rect 4895 19552 4911 19616
rect 4975 19552 4991 19616
rect 5055 19552 5071 19616
rect 5135 19552 5141 19616
rect 4825 19551 5141 19552
rect 11264 19616 11580 19617
rect 11264 19552 11270 19616
rect 11334 19552 11350 19616
rect 11414 19552 11430 19616
rect 11494 19552 11510 19616
rect 11574 19552 11580 19616
rect 11264 19551 11580 19552
rect 17703 19616 18019 19617
rect 17703 19552 17709 19616
rect 17773 19552 17789 19616
rect 17853 19552 17869 19616
rect 17933 19552 17949 19616
rect 18013 19552 18019 19616
rect 17703 19551 18019 19552
rect 24142 19616 24458 19617
rect 24142 19552 24148 19616
rect 24212 19552 24228 19616
rect 24292 19552 24308 19616
rect 24372 19552 24388 19616
rect 24452 19552 24458 19616
rect 24142 19551 24458 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 5257 19410 5323 19413
rect 10409 19410 10475 19413
rect 5257 19408 10475 19410
rect 5257 19352 5262 19408
rect 5318 19352 10414 19408
rect 10470 19352 10475 19408
rect 5257 19350 10475 19352
rect 5257 19347 5323 19350
rect 10409 19347 10475 19350
rect 4165 19072 4481 19073
rect 4165 19008 4171 19072
rect 4235 19008 4251 19072
rect 4315 19008 4331 19072
rect 4395 19008 4411 19072
rect 4475 19008 4481 19072
rect 4165 19007 4481 19008
rect 10604 19072 10920 19073
rect 10604 19008 10610 19072
rect 10674 19008 10690 19072
rect 10754 19008 10770 19072
rect 10834 19008 10850 19072
rect 10914 19008 10920 19072
rect 10604 19007 10920 19008
rect 17043 19072 17359 19073
rect 17043 19008 17049 19072
rect 17113 19008 17129 19072
rect 17193 19008 17209 19072
rect 17273 19008 17289 19072
rect 17353 19008 17359 19072
rect 17043 19007 17359 19008
rect 23482 19072 23798 19073
rect 23482 19008 23488 19072
rect 23552 19008 23568 19072
rect 23632 19008 23648 19072
rect 23712 19008 23728 19072
rect 23792 19008 23798 19072
rect 23482 19007 23798 19008
rect 15101 18866 15167 18869
rect 17953 18866 18019 18869
rect 15101 18864 18019 18866
rect 15101 18808 15106 18864
rect 15162 18808 17958 18864
rect 18014 18808 18019 18864
rect 15101 18806 18019 18808
rect 15101 18803 15167 18806
rect 17953 18803 18019 18806
rect 26509 18594 26575 18597
rect 27188 18594 27988 18624
rect 26509 18592 27988 18594
rect 26509 18536 26514 18592
rect 26570 18536 27988 18592
rect 26509 18534 27988 18536
rect 26509 18531 26575 18534
rect 4825 18528 5141 18529
rect 4825 18464 4831 18528
rect 4895 18464 4911 18528
rect 4975 18464 4991 18528
rect 5055 18464 5071 18528
rect 5135 18464 5141 18528
rect 4825 18463 5141 18464
rect 11264 18528 11580 18529
rect 11264 18464 11270 18528
rect 11334 18464 11350 18528
rect 11414 18464 11430 18528
rect 11494 18464 11510 18528
rect 11574 18464 11580 18528
rect 11264 18463 11580 18464
rect 17703 18528 18019 18529
rect 17703 18464 17709 18528
rect 17773 18464 17789 18528
rect 17853 18464 17869 18528
rect 17933 18464 17949 18528
rect 18013 18464 18019 18528
rect 17703 18463 18019 18464
rect 24142 18528 24458 18529
rect 24142 18464 24148 18528
rect 24212 18464 24228 18528
rect 24292 18464 24308 18528
rect 24372 18464 24388 18528
rect 24452 18464 24458 18528
rect 27188 18504 27988 18534
rect 24142 18463 24458 18464
rect 4165 17984 4481 17985
rect 4165 17920 4171 17984
rect 4235 17920 4251 17984
rect 4315 17920 4331 17984
rect 4395 17920 4411 17984
rect 4475 17920 4481 17984
rect 4165 17919 4481 17920
rect 10604 17984 10920 17985
rect 10604 17920 10610 17984
rect 10674 17920 10690 17984
rect 10754 17920 10770 17984
rect 10834 17920 10850 17984
rect 10914 17920 10920 17984
rect 10604 17919 10920 17920
rect 17043 17984 17359 17985
rect 17043 17920 17049 17984
rect 17113 17920 17129 17984
rect 17193 17920 17209 17984
rect 17273 17920 17289 17984
rect 17353 17920 17359 17984
rect 17043 17919 17359 17920
rect 23482 17984 23798 17985
rect 23482 17920 23488 17984
rect 23552 17920 23568 17984
rect 23632 17920 23648 17984
rect 23712 17920 23728 17984
rect 23792 17920 23798 17984
rect 23482 17919 23798 17920
rect 15469 17916 15535 17917
rect 15469 17914 15516 17916
rect 15424 17912 15516 17914
rect 15424 17856 15474 17912
rect 15424 17854 15516 17856
rect 15469 17852 15516 17854
rect 15580 17852 15586 17916
rect 15469 17851 15535 17852
rect 4825 17440 5141 17441
rect 4825 17376 4831 17440
rect 4895 17376 4911 17440
rect 4975 17376 4991 17440
rect 5055 17376 5071 17440
rect 5135 17376 5141 17440
rect 4825 17375 5141 17376
rect 11264 17440 11580 17441
rect 11264 17376 11270 17440
rect 11334 17376 11350 17440
rect 11414 17376 11430 17440
rect 11494 17376 11510 17440
rect 11574 17376 11580 17440
rect 11264 17375 11580 17376
rect 17703 17440 18019 17441
rect 17703 17376 17709 17440
rect 17773 17376 17789 17440
rect 17853 17376 17869 17440
rect 17933 17376 17949 17440
rect 18013 17376 18019 17440
rect 17703 17375 18019 17376
rect 24142 17440 24458 17441
rect 24142 17376 24148 17440
rect 24212 17376 24228 17440
rect 24292 17376 24308 17440
rect 24372 17376 24388 17440
rect 24452 17376 24458 17440
rect 24142 17375 24458 17376
rect 15377 17372 15443 17373
rect 15326 17308 15332 17372
rect 15396 17370 15443 17372
rect 15396 17368 15488 17370
rect 15438 17312 15488 17368
rect 15396 17310 15488 17312
rect 15396 17308 15443 17310
rect 15377 17307 15443 17308
rect 0 17234 800 17264
rect 933 17234 999 17237
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 0 17144 800 17174
rect 933 17171 999 17174
rect 13169 17234 13235 17237
rect 18781 17234 18847 17237
rect 13169 17232 18847 17234
rect 13169 17176 13174 17232
rect 13230 17176 18786 17232
rect 18842 17176 18847 17232
rect 13169 17174 18847 17176
rect 13169 17171 13235 17174
rect 18781 17171 18847 17174
rect 4165 16896 4481 16897
rect 4165 16832 4171 16896
rect 4235 16832 4251 16896
rect 4315 16832 4331 16896
rect 4395 16832 4411 16896
rect 4475 16832 4481 16896
rect 4165 16831 4481 16832
rect 10604 16896 10920 16897
rect 10604 16832 10610 16896
rect 10674 16832 10690 16896
rect 10754 16832 10770 16896
rect 10834 16832 10850 16896
rect 10914 16832 10920 16896
rect 10604 16831 10920 16832
rect 17043 16896 17359 16897
rect 17043 16832 17049 16896
rect 17113 16832 17129 16896
rect 17193 16832 17209 16896
rect 17273 16832 17289 16896
rect 17353 16832 17359 16896
rect 17043 16831 17359 16832
rect 23482 16896 23798 16897
rect 23482 16832 23488 16896
rect 23552 16832 23568 16896
rect 23632 16832 23648 16896
rect 23712 16832 23728 16896
rect 23792 16832 23798 16896
rect 23482 16831 23798 16832
rect 4825 16352 5141 16353
rect 4825 16288 4831 16352
rect 4895 16288 4911 16352
rect 4975 16288 4991 16352
rect 5055 16288 5071 16352
rect 5135 16288 5141 16352
rect 4825 16287 5141 16288
rect 11264 16352 11580 16353
rect 11264 16288 11270 16352
rect 11334 16288 11350 16352
rect 11414 16288 11430 16352
rect 11494 16288 11510 16352
rect 11574 16288 11580 16352
rect 11264 16287 11580 16288
rect 17703 16352 18019 16353
rect 17703 16288 17709 16352
rect 17773 16288 17789 16352
rect 17853 16288 17869 16352
rect 17933 16288 17949 16352
rect 18013 16288 18019 16352
rect 17703 16287 18019 16288
rect 24142 16352 24458 16353
rect 24142 16288 24148 16352
rect 24212 16288 24228 16352
rect 24292 16288 24308 16352
rect 24372 16288 24388 16352
rect 24452 16288 24458 16352
rect 24142 16287 24458 16288
rect 11329 16146 11395 16149
rect 13169 16146 13235 16149
rect 11329 16144 13235 16146
rect 11329 16088 11334 16144
rect 11390 16088 13174 16144
rect 13230 16088 13235 16144
rect 11329 16086 13235 16088
rect 11329 16083 11395 16086
rect 13169 16083 13235 16086
rect 17401 16146 17467 16149
rect 17677 16146 17743 16149
rect 18413 16146 18479 16149
rect 17401 16144 18479 16146
rect 17401 16088 17406 16144
rect 17462 16088 17682 16144
rect 17738 16088 18418 16144
rect 18474 16088 18479 16144
rect 17401 16086 18479 16088
rect 17401 16083 17467 16086
rect 17677 16083 17743 16086
rect 18413 16083 18479 16086
rect 1577 16010 1643 16013
rect 7373 16010 7439 16013
rect 1577 16008 7439 16010
rect 1577 15952 1582 16008
rect 1638 15952 7378 16008
rect 7434 15952 7439 16008
rect 1577 15950 7439 15952
rect 1577 15947 1643 15950
rect 7373 15947 7439 15950
rect 4165 15808 4481 15809
rect 4165 15744 4171 15808
rect 4235 15744 4251 15808
rect 4315 15744 4331 15808
rect 4395 15744 4411 15808
rect 4475 15744 4481 15808
rect 4165 15743 4481 15744
rect 10604 15808 10920 15809
rect 10604 15744 10610 15808
rect 10674 15744 10690 15808
rect 10754 15744 10770 15808
rect 10834 15744 10850 15808
rect 10914 15744 10920 15808
rect 10604 15743 10920 15744
rect 17043 15808 17359 15809
rect 17043 15744 17049 15808
rect 17113 15744 17129 15808
rect 17193 15744 17209 15808
rect 17273 15744 17289 15808
rect 17353 15744 17359 15808
rect 17043 15743 17359 15744
rect 23482 15808 23798 15809
rect 23482 15744 23488 15808
rect 23552 15744 23568 15808
rect 23632 15744 23648 15808
rect 23712 15744 23728 15808
rect 23792 15744 23798 15808
rect 23482 15743 23798 15744
rect 4825 15264 5141 15265
rect 4825 15200 4831 15264
rect 4895 15200 4911 15264
rect 4975 15200 4991 15264
rect 5055 15200 5071 15264
rect 5135 15200 5141 15264
rect 4825 15199 5141 15200
rect 11264 15264 11580 15265
rect 11264 15200 11270 15264
rect 11334 15200 11350 15264
rect 11414 15200 11430 15264
rect 11494 15200 11510 15264
rect 11574 15200 11580 15264
rect 11264 15199 11580 15200
rect 17703 15264 18019 15265
rect 17703 15200 17709 15264
rect 17773 15200 17789 15264
rect 17853 15200 17869 15264
rect 17933 15200 17949 15264
rect 18013 15200 18019 15264
rect 17703 15199 18019 15200
rect 24142 15264 24458 15265
rect 24142 15200 24148 15264
rect 24212 15200 24228 15264
rect 24292 15200 24308 15264
rect 24372 15200 24388 15264
rect 24452 15200 24458 15264
rect 24142 15199 24458 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 4165 14720 4481 14721
rect 4165 14656 4171 14720
rect 4235 14656 4251 14720
rect 4315 14656 4331 14720
rect 4395 14656 4411 14720
rect 4475 14656 4481 14720
rect 4165 14655 4481 14656
rect 10604 14720 10920 14721
rect 10604 14656 10610 14720
rect 10674 14656 10690 14720
rect 10754 14656 10770 14720
rect 10834 14656 10850 14720
rect 10914 14656 10920 14720
rect 10604 14655 10920 14656
rect 17043 14720 17359 14721
rect 17043 14656 17049 14720
rect 17113 14656 17129 14720
rect 17193 14656 17209 14720
rect 17273 14656 17289 14720
rect 17353 14656 17359 14720
rect 17043 14655 17359 14656
rect 23482 14720 23798 14721
rect 23482 14656 23488 14720
rect 23552 14656 23568 14720
rect 23632 14656 23648 14720
rect 23712 14656 23728 14720
rect 23792 14656 23798 14720
rect 23482 14655 23798 14656
rect 17217 14514 17283 14517
rect 17953 14514 18019 14517
rect 17217 14512 18019 14514
rect 17217 14456 17222 14512
rect 17278 14456 17958 14512
rect 18014 14456 18019 14512
rect 17217 14454 18019 14456
rect 17217 14451 17283 14454
rect 17953 14451 18019 14454
rect 18321 14514 18387 14517
rect 19057 14514 19123 14517
rect 18321 14512 19123 14514
rect 18321 14456 18326 14512
rect 18382 14456 19062 14512
rect 19118 14456 19123 14512
rect 18321 14454 19123 14456
rect 18321 14451 18387 14454
rect 19057 14451 19123 14454
rect 15653 14378 15719 14381
rect 18781 14378 18847 14381
rect 15653 14376 18847 14378
rect 15653 14320 15658 14376
rect 15714 14320 18786 14376
rect 18842 14320 18847 14376
rect 15653 14318 18847 14320
rect 15653 14315 15719 14318
rect 18781 14315 18847 14318
rect 4825 14176 5141 14177
rect 4825 14112 4831 14176
rect 4895 14112 4911 14176
rect 4975 14112 4991 14176
rect 5055 14112 5071 14176
rect 5135 14112 5141 14176
rect 4825 14111 5141 14112
rect 11264 14176 11580 14177
rect 11264 14112 11270 14176
rect 11334 14112 11350 14176
rect 11414 14112 11430 14176
rect 11494 14112 11510 14176
rect 11574 14112 11580 14176
rect 11264 14111 11580 14112
rect 17703 14176 18019 14177
rect 17703 14112 17709 14176
rect 17773 14112 17789 14176
rect 17853 14112 17869 14176
rect 17933 14112 17949 14176
rect 18013 14112 18019 14176
rect 17703 14111 18019 14112
rect 24142 14176 24458 14177
rect 24142 14112 24148 14176
rect 24212 14112 24228 14176
rect 24292 14112 24308 14176
rect 24372 14112 24388 14176
rect 24452 14112 24458 14176
rect 24142 14111 24458 14112
rect 4165 13632 4481 13633
rect 4165 13568 4171 13632
rect 4235 13568 4251 13632
rect 4315 13568 4331 13632
rect 4395 13568 4411 13632
rect 4475 13568 4481 13632
rect 4165 13567 4481 13568
rect 10604 13632 10920 13633
rect 10604 13568 10610 13632
rect 10674 13568 10690 13632
rect 10754 13568 10770 13632
rect 10834 13568 10850 13632
rect 10914 13568 10920 13632
rect 10604 13567 10920 13568
rect 17043 13632 17359 13633
rect 17043 13568 17049 13632
rect 17113 13568 17129 13632
rect 17193 13568 17209 13632
rect 17273 13568 17289 13632
rect 17353 13568 17359 13632
rect 17043 13567 17359 13568
rect 23482 13632 23798 13633
rect 23482 13568 23488 13632
rect 23552 13568 23568 13632
rect 23632 13568 23648 13632
rect 23712 13568 23728 13632
rect 23792 13568 23798 13632
rect 23482 13567 23798 13568
rect 7649 13426 7715 13429
rect 12525 13426 12591 13429
rect 7649 13424 12591 13426
rect 7649 13368 7654 13424
rect 7710 13368 12530 13424
rect 12586 13368 12591 13424
rect 7649 13366 12591 13368
rect 7649 13363 7715 13366
rect 12525 13363 12591 13366
rect 5073 13290 5139 13293
rect 8845 13290 8911 13293
rect 5073 13288 8911 13290
rect 5073 13232 5078 13288
rect 5134 13232 8850 13288
rect 8906 13232 8911 13288
rect 5073 13230 8911 13232
rect 5073 13227 5139 13230
rect 8845 13227 8911 13230
rect 9029 13290 9095 13293
rect 9305 13290 9371 13293
rect 20989 13290 21055 13293
rect 9029 13288 21055 13290
rect 9029 13232 9034 13288
rect 9090 13232 9310 13288
rect 9366 13232 20994 13288
rect 21050 13232 21055 13288
rect 9029 13230 21055 13232
rect 9029 13227 9095 13230
rect 9305 13227 9371 13230
rect 20989 13227 21055 13230
rect 4825 13088 5141 13089
rect 4825 13024 4831 13088
rect 4895 13024 4911 13088
rect 4975 13024 4991 13088
rect 5055 13024 5071 13088
rect 5135 13024 5141 13088
rect 4825 13023 5141 13024
rect 11264 13088 11580 13089
rect 11264 13024 11270 13088
rect 11334 13024 11350 13088
rect 11414 13024 11430 13088
rect 11494 13024 11510 13088
rect 11574 13024 11580 13088
rect 11264 13023 11580 13024
rect 17703 13088 18019 13089
rect 17703 13024 17709 13088
rect 17773 13024 17789 13088
rect 17853 13024 17869 13088
rect 17933 13024 17949 13088
rect 18013 13024 18019 13088
rect 17703 13023 18019 13024
rect 24142 13088 24458 13089
rect 24142 13024 24148 13088
rect 24212 13024 24228 13088
rect 24292 13024 24308 13088
rect 24372 13024 24388 13088
rect 24452 13024 24458 13088
rect 24142 13023 24458 13024
rect 0 12882 800 12912
rect 1393 12882 1459 12885
rect 0 12880 1459 12882
rect 0 12824 1398 12880
rect 1454 12824 1459 12880
rect 0 12822 1459 12824
rect 0 12792 800 12822
rect 1393 12819 1459 12822
rect 3969 12882 4035 12885
rect 13077 12882 13143 12885
rect 3969 12880 13143 12882
rect 3969 12824 3974 12880
rect 4030 12824 13082 12880
rect 13138 12824 13143 12880
rect 3969 12822 13143 12824
rect 3969 12819 4035 12822
rect 13077 12819 13143 12822
rect 8845 12746 8911 12749
rect 14457 12746 14523 12749
rect 15101 12746 15167 12749
rect 8845 12744 15167 12746
rect 8845 12688 8850 12744
rect 8906 12688 14462 12744
rect 14518 12688 15106 12744
rect 15162 12688 15167 12744
rect 8845 12686 15167 12688
rect 8845 12683 8911 12686
rect 14457 12683 14523 12686
rect 15101 12683 15167 12686
rect 4165 12544 4481 12545
rect 4165 12480 4171 12544
rect 4235 12480 4251 12544
rect 4315 12480 4331 12544
rect 4395 12480 4411 12544
rect 4475 12480 4481 12544
rect 4165 12479 4481 12480
rect 10604 12544 10920 12545
rect 10604 12480 10610 12544
rect 10674 12480 10690 12544
rect 10754 12480 10770 12544
rect 10834 12480 10850 12544
rect 10914 12480 10920 12544
rect 10604 12479 10920 12480
rect 17043 12544 17359 12545
rect 17043 12480 17049 12544
rect 17113 12480 17129 12544
rect 17193 12480 17209 12544
rect 17273 12480 17289 12544
rect 17353 12480 17359 12544
rect 17043 12479 17359 12480
rect 23482 12544 23798 12545
rect 23482 12480 23488 12544
rect 23552 12480 23568 12544
rect 23632 12480 23648 12544
rect 23712 12480 23728 12544
rect 23792 12480 23798 12544
rect 23482 12479 23798 12480
rect 4825 12000 5141 12001
rect 4825 11936 4831 12000
rect 4895 11936 4911 12000
rect 4975 11936 4991 12000
rect 5055 11936 5071 12000
rect 5135 11936 5141 12000
rect 4825 11935 5141 11936
rect 11264 12000 11580 12001
rect 11264 11936 11270 12000
rect 11334 11936 11350 12000
rect 11414 11936 11430 12000
rect 11494 11936 11510 12000
rect 11574 11936 11580 12000
rect 11264 11935 11580 11936
rect 17703 12000 18019 12001
rect 17703 11936 17709 12000
rect 17773 11936 17789 12000
rect 17853 11936 17869 12000
rect 17933 11936 17949 12000
rect 18013 11936 18019 12000
rect 17703 11935 18019 11936
rect 24142 12000 24458 12001
rect 24142 11936 24148 12000
rect 24212 11936 24228 12000
rect 24292 11936 24308 12000
rect 24372 11936 24388 12000
rect 24452 11936 24458 12000
rect 24142 11935 24458 11936
rect 15193 11794 15259 11797
rect 16849 11794 16915 11797
rect 18781 11794 18847 11797
rect 15193 11792 18847 11794
rect 15193 11736 15198 11792
rect 15254 11736 16854 11792
rect 16910 11736 18786 11792
rect 18842 11736 18847 11792
rect 15193 11734 18847 11736
rect 15193 11731 15259 11734
rect 16849 11731 16915 11734
rect 18781 11731 18847 11734
rect 4165 11456 4481 11457
rect 4165 11392 4171 11456
rect 4235 11392 4251 11456
rect 4315 11392 4331 11456
rect 4395 11392 4411 11456
rect 4475 11392 4481 11456
rect 4165 11391 4481 11392
rect 10604 11456 10920 11457
rect 10604 11392 10610 11456
rect 10674 11392 10690 11456
rect 10754 11392 10770 11456
rect 10834 11392 10850 11456
rect 10914 11392 10920 11456
rect 10604 11391 10920 11392
rect 17043 11456 17359 11457
rect 17043 11392 17049 11456
rect 17113 11392 17129 11456
rect 17193 11392 17209 11456
rect 17273 11392 17289 11456
rect 17353 11392 17359 11456
rect 17043 11391 17359 11392
rect 23482 11456 23798 11457
rect 23482 11392 23488 11456
rect 23552 11392 23568 11456
rect 23632 11392 23648 11456
rect 23712 11392 23728 11456
rect 23792 11392 23798 11456
rect 23482 11391 23798 11392
rect 26509 11250 26575 11253
rect 27188 11250 27988 11280
rect 26509 11248 27988 11250
rect 26509 11192 26514 11248
rect 26570 11192 27988 11248
rect 26509 11190 27988 11192
rect 26509 11187 26575 11190
rect 27188 11160 27988 11190
rect 4061 11114 4127 11117
rect 6729 11114 6795 11117
rect 4061 11112 6795 11114
rect 4061 11056 4066 11112
rect 4122 11056 6734 11112
rect 6790 11056 6795 11112
rect 4061 11054 6795 11056
rect 4061 11051 4127 11054
rect 6729 11051 6795 11054
rect 4825 10912 5141 10913
rect 4825 10848 4831 10912
rect 4895 10848 4911 10912
rect 4975 10848 4991 10912
rect 5055 10848 5071 10912
rect 5135 10848 5141 10912
rect 4825 10847 5141 10848
rect 11264 10912 11580 10913
rect 11264 10848 11270 10912
rect 11334 10848 11350 10912
rect 11414 10848 11430 10912
rect 11494 10848 11510 10912
rect 11574 10848 11580 10912
rect 11264 10847 11580 10848
rect 17703 10912 18019 10913
rect 17703 10848 17709 10912
rect 17773 10848 17789 10912
rect 17853 10848 17869 10912
rect 17933 10848 17949 10912
rect 18013 10848 18019 10912
rect 17703 10847 18019 10848
rect 24142 10912 24458 10913
rect 24142 10848 24148 10912
rect 24212 10848 24228 10912
rect 24292 10848 24308 10912
rect 24372 10848 24388 10912
rect 24452 10848 24458 10912
rect 24142 10847 24458 10848
rect 0 10706 800 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 800 10646
rect 1393 10643 1459 10646
rect 4165 10368 4481 10369
rect 4165 10304 4171 10368
rect 4235 10304 4251 10368
rect 4315 10304 4331 10368
rect 4395 10304 4411 10368
rect 4475 10304 4481 10368
rect 4165 10303 4481 10304
rect 10604 10368 10920 10369
rect 10604 10304 10610 10368
rect 10674 10304 10690 10368
rect 10754 10304 10770 10368
rect 10834 10304 10850 10368
rect 10914 10304 10920 10368
rect 10604 10303 10920 10304
rect 17043 10368 17359 10369
rect 17043 10304 17049 10368
rect 17113 10304 17129 10368
rect 17193 10304 17209 10368
rect 17273 10304 17289 10368
rect 17353 10304 17359 10368
rect 17043 10303 17359 10304
rect 23482 10368 23798 10369
rect 23482 10304 23488 10368
rect 23552 10304 23568 10368
rect 23632 10304 23648 10368
rect 23712 10304 23728 10368
rect 23792 10304 23798 10368
rect 23482 10303 23798 10304
rect 4797 10026 4863 10029
rect 5349 10026 5415 10029
rect 4797 10024 5415 10026
rect 4797 9968 4802 10024
rect 4858 9968 5354 10024
rect 5410 9968 5415 10024
rect 4797 9966 5415 9968
rect 4797 9963 4863 9966
rect 5349 9963 5415 9966
rect 4825 9824 5141 9825
rect 4825 9760 4831 9824
rect 4895 9760 4911 9824
rect 4975 9760 4991 9824
rect 5055 9760 5071 9824
rect 5135 9760 5141 9824
rect 4825 9759 5141 9760
rect 11264 9824 11580 9825
rect 11264 9760 11270 9824
rect 11334 9760 11350 9824
rect 11414 9760 11430 9824
rect 11494 9760 11510 9824
rect 11574 9760 11580 9824
rect 11264 9759 11580 9760
rect 17703 9824 18019 9825
rect 17703 9760 17709 9824
rect 17773 9760 17789 9824
rect 17853 9760 17869 9824
rect 17933 9760 17949 9824
rect 18013 9760 18019 9824
rect 17703 9759 18019 9760
rect 24142 9824 24458 9825
rect 24142 9760 24148 9824
rect 24212 9760 24228 9824
rect 24292 9760 24308 9824
rect 24372 9760 24388 9824
rect 24452 9760 24458 9824
rect 24142 9759 24458 9760
rect 4165 9280 4481 9281
rect 4165 9216 4171 9280
rect 4235 9216 4251 9280
rect 4315 9216 4331 9280
rect 4395 9216 4411 9280
rect 4475 9216 4481 9280
rect 4165 9215 4481 9216
rect 10604 9280 10920 9281
rect 10604 9216 10610 9280
rect 10674 9216 10690 9280
rect 10754 9216 10770 9280
rect 10834 9216 10850 9280
rect 10914 9216 10920 9280
rect 10604 9215 10920 9216
rect 17043 9280 17359 9281
rect 17043 9216 17049 9280
rect 17113 9216 17129 9280
rect 17193 9216 17209 9280
rect 17273 9216 17289 9280
rect 17353 9216 17359 9280
rect 17043 9215 17359 9216
rect 23482 9280 23798 9281
rect 23482 9216 23488 9280
rect 23552 9216 23568 9280
rect 23632 9216 23648 9280
rect 23712 9216 23728 9280
rect 23792 9216 23798 9280
rect 23482 9215 23798 9216
rect 11053 9210 11119 9213
rect 12985 9210 13051 9213
rect 11053 9208 13051 9210
rect 11053 9152 11058 9208
rect 11114 9152 12990 9208
rect 13046 9152 13051 9208
rect 11053 9150 13051 9152
rect 11053 9147 11119 9150
rect 12985 9147 13051 9150
rect 10777 8938 10843 8941
rect 13261 8938 13327 8941
rect 10777 8936 13327 8938
rect 10777 8880 10782 8936
rect 10838 8880 13266 8936
rect 13322 8880 13327 8936
rect 10777 8878 13327 8880
rect 10777 8875 10843 8878
rect 13261 8875 13327 8878
rect 4825 8736 5141 8737
rect 4825 8672 4831 8736
rect 4895 8672 4911 8736
rect 4975 8672 4991 8736
rect 5055 8672 5071 8736
rect 5135 8672 5141 8736
rect 4825 8671 5141 8672
rect 11264 8736 11580 8737
rect 11264 8672 11270 8736
rect 11334 8672 11350 8736
rect 11414 8672 11430 8736
rect 11494 8672 11510 8736
rect 11574 8672 11580 8736
rect 11264 8671 11580 8672
rect 17703 8736 18019 8737
rect 17703 8672 17709 8736
rect 17773 8672 17789 8736
rect 17853 8672 17869 8736
rect 17933 8672 17949 8736
rect 18013 8672 18019 8736
rect 17703 8671 18019 8672
rect 24142 8736 24458 8737
rect 24142 8672 24148 8736
rect 24212 8672 24228 8736
rect 24292 8672 24308 8736
rect 24372 8672 24388 8736
rect 24452 8672 24458 8736
rect 24142 8671 24458 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 4165 8192 4481 8193
rect 4165 8128 4171 8192
rect 4235 8128 4251 8192
rect 4315 8128 4331 8192
rect 4395 8128 4411 8192
rect 4475 8128 4481 8192
rect 4165 8127 4481 8128
rect 10604 8192 10920 8193
rect 10604 8128 10610 8192
rect 10674 8128 10690 8192
rect 10754 8128 10770 8192
rect 10834 8128 10850 8192
rect 10914 8128 10920 8192
rect 10604 8127 10920 8128
rect 17043 8192 17359 8193
rect 17043 8128 17049 8192
rect 17113 8128 17129 8192
rect 17193 8128 17209 8192
rect 17273 8128 17289 8192
rect 17353 8128 17359 8192
rect 17043 8127 17359 8128
rect 23482 8192 23798 8193
rect 23482 8128 23488 8192
rect 23552 8128 23568 8192
rect 23632 8128 23648 8192
rect 23712 8128 23728 8192
rect 23792 8128 23798 8192
rect 23482 8127 23798 8128
rect 4825 7648 5141 7649
rect 4825 7584 4831 7648
rect 4895 7584 4911 7648
rect 4975 7584 4991 7648
rect 5055 7584 5071 7648
rect 5135 7584 5141 7648
rect 4825 7583 5141 7584
rect 11264 7648 11580 7649
rect 11264 7584 11270 7648
rect 11334 7584 11350 7648
rect 11414 7584 11430 7648
rect 11494 7584 11510 7648
rect 11574 7584 11580 7648
rect 11264 7583 11580 7584
rect 17703 7648 18019 7649
rect 17703 7584 17709 7648
rect 17773 7584 17789 7648
rect 17853 7584 17869 7648
rect 17933 7584 17949 7648
rect 18013 7584 18019 7648
rect 17703 7583 18019 7584
rect 24142 7648 24458 7649
rect 24142 7584 24148 7648
rect 24212 7584 24228 7648
rect 24292 7584 24308 7648
rect 24372 7584 24388 7648
rect 24452 7584 24458 7648
rect 24142 7583 24458 7584
rect 11789 7442 11855 7445
rect 25681 7442 25747 7445
rect 11789 7440 25747 7442
rect 11789 7384 11794 7440
rect 11850 7384 25686 7440
rect 25742 7384 25747 7440
rect 11789 7382 25747 7384
rect 11789 7379 11855 7382
rect 25681 7379 25747 7382
rect 9121 7306 9187 7309
rect 10317 7306 10383 7309
rect 9121 7304 10383 7306
rect 9121 7248 9126 7304
rect 9182 7248 10322 7304
rect 10378 7248 10383 7304
rect 9121 7246 10383 7248
rect 9121 7243 9187 7246
rect 10317 7243 10383 7246
rect 10593 7306 10659 7309
rect 17033 7306 17099 7309
rect 10593 7304 17099 7306
rect 10593 7248 10598 7304
rect 10654 7248 17038 7304
rect 17094 7248 17099 7304
rect 10593 7246 17099 7248
rect 10593 7243 10659 7246
rect 17033 7243 17099 7246
rect 4165 7104 4481 7105
rect 4165 7040 4171 7104
rect 4235 7040 4251 7104
rect 4315 7040 4331 7104
rect 4395 7040 4411 7104
rect 4475 7040 4481 7104
rect 4165 7039 4481 7040
rect 10604 7104 10920 7105
rect 10604 7040 10610 7104
rect 10674 7040 10690 7104
rect 10754 7040 10770 7104
rect 10834 7040 10850 7104
rect 10914 7040 10920 7104
rect 10604 7039 10920 7040
rect 17043 7104 17359 7105
rect 17043 7040 17049 7104
rect 17113 7040 17129 7104
rect 17193 7040 17209 7104
rect 17273 7040 17289 7104
rect 17353 7040 17359 7104
rect 17043 7039 17359 7040
rect 23482 7104 23798 7105
rect 23482 7040 23488 7104
rect 23552 7040 23568 7104
rect 23632 7040 23648 7104
rect 23712 7040 23728 7104
rect 23792 7040 23798 7104
rect 23482 7039 23798 7040
rect 9581 6898 9647 6901
rect 14365 6898 14431 6901
rect 9581 6896 14431 6898
rect 9581 6840 9586 6896
rect 9642 6840 14370 6896
rect 14426 6840 14431 6896
rect 9581 6838 14431 6840
rect 9581 6835 9647 6838
rect 14365 6835 14431 6838
rect 8477 6762 8543 6765
rect 15193 6762 15259 6765
rect 8477 6760 15259 6762
rect 8477 6704 8482 6760
rect 8538 6704 15198 6760
rect 15254 6704 15259 6760
rect 8477 6702 15259 6704
rect 8477 6699 8543 6702
rect 15193 6699 15259 6702
rect 9673 6626 9739 6629
rect 10225 6626 10291 6629
rect 9673 6624 10291 6626
rect 9673 6568 9678 6624
rect 9734 6568 10230 6624
rect 10286 6568 10291 6624
rect 9673 6566 10291 6568
rect 9673 6563 9739 6566
rect 10225 6563 10291 6566
rect 4825 6560 5141 6561
rect 4825 6496 4831 6560
rect 4895 6496 4911 6560
rect 4975 6496 4991 6560
rect 5055 6496 5071 6560
rect 5135 6496 5141 6560
rect 4825 6495 5141 6496
rect 11264 6560 11580 6561
rect 11264 6496 11270 6560
rect 11334 6496 11350 6560
rect 11414 6496 11430 6560
rect 11494 6496 11510 6560
rect 11574 6496 11580 6560
rect 11264 6495 11580 6496
rect 17703 6560 18019 6561
rect 17703 6496 17709 6560
rect 17773 6496 17789 6560
rect 17853 6496 17869 6560
rect 17933 6496 17949 6560
rect 18013 6496 18019 6560
rect 17703 6495 18019 6496
rect 24142 6560 24458 6561
rect 24142 6496 24148 6560
rect 24212 6496 24228 6560
rect 24292 6496 24308 6560
rect 24372 6496 24388 6560
rect 24452 6496 24458 6560
rect 24142 6495 24458 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 8937 6354 9003 6357
rect 9949 6354 10015 6357
rect 8937 6352 10015 6354
rect 8937 6296 8942 6352
rect 8998 6296 9954 6352
rect 10010 6296 10015 6352
rect 8937 6294 10015 6296
rect 8937 6291 9003 6294
rect 9949 6291 10015 6294
rect 4165 6016 4481 6017
rect 4165 5952 4171 6016
rect 4235 5952 4251 6016
rect 4315 5952 4331 6016
rect 4395 5952 4411 6016
rect 4475 5952 4481 6016
rect 4165 5951 4481 5952
rect 10604 6016 10920 6017
rect 10604 5952 10610 6016
rect 10674 5952 10690 6016
rect 10754 5952 10770 6016
rect 10834 5952 10850 6016
rect 10914 5952 10920 6016
rect 10604 5951 10920 5952
rect 17043 6016 17359 6017
rect 17043 5952 17049 6016
rect 17113 5952 17129 6016
rect 17193 5952 17209 6016
rect 17273 5952 17289 6016
rect 17353 5952 17359 6016
rect 17043 5951 17359 5952
rect 23482 6016 23798 6017
rect 23482 5952 23488 6016
rect 23552 5952 23568 6016
rect 23632 5952 23648 6016
rect 23712 5952 23728 6016
rect 23792 5952 23798 6016
rect 23482 5951 23798 5952
rect 4825 5472 5141 5473
rect 4825 5408 4831 5472
rect 4895 5408 4911 5472
rect 4975 5408 4991 5472
rect 5055 5408 5071 5472
rect 5135 5408 5141 5472
rect 4825 5407 5141 5408
rect 11264 5472 11580 5473
rect 11264 5408 11270 5472
rect 11334 5408 11350 5472
rect 11414 5408 11430 5472
rect 11494 5408 11510 5472
rect 11574 5408 11580 5472
rect 11264 5407 11580 5408
rect 17703 5472 18019 5473
rect 17703 5408 17709 5472
rect 17773 5408 17789 5472
rect 17853 5408 17869 5472
rect 17933 5408 17949 5472
rect 18013 5408 18019 5472
rect 17703 5407 18019 5408
rect 24142 5472 24458 5473
rect 24142 5408 24148 5472
rect 24212 5408 24228 5472
rect 24292 5408 24308 5472
rect 24372 5408 24388 5472
rect 24452 5408 24458 5472
rect 24142 5407 24458 5408
rect 13629 5266 13695 5269
rect 15101 5266 15167 5269
rect 13629 5264 15167 5266
rect 13629 5208 13634 5264
rect 13690 5208 15106 5264
rect 15162 5208 15167 5264
rect 13629 5206 15167 5208
rect 13629 5203 13695 5206
rect 15101 5203 15167 5206
rect 4165 4928 4481 4929
rect 4165 4864 4171 4928
rect 4235 4864 4251 4928
rect 4315 4864 4331 4928
rect 4395 4864 4411 4928
rect 4475 4864 4481 4928
rect 4165 4863 4481 4864
rect 10604 4928 10920 4929
rect 10604 4864 10610 4928
rect 10674 4864 10690 4928
rect 10754 4864 10770 4928
rect 10834 4864 10850 4928
rect 10914 4864 10920 4928
rect 10604 4863 10920 4864
rect 17043 4928 17359 4929
rect 17043 4864 17049 4928
rect 17113 4864 17129 4928
rect 17193 4864 17209 4928
rect 17273 4864 17289 4928
rect 17353 4864 17359 4928
rect 17043 4863 17359 4864
rect 23482 4928 23798 4929
rect 23482 4864 23488 4928
rect 23552 4864 23568 4928
rect 23632 4864 23648 4928
rect 23712 4864 23728 4928
rect 23792 4864 23798 4928
rect 23482 4863 23798 4864
rect 11053 4586 11119 4589
rect 13077 4586 13143 4589
rect 11053 4584 13143 4586
rect 11053 4528 11058 4584
rect 11114 4528 13082 4584
rect 13138 4528 13143 4584
rect 11053 4526 13143 4528
rect 11053 4523 11119 4526
rect 13077 4523 13143 4526
rect 14365 4450 14431 4453
rect 16757 4450 16823 4453
rect 14365 4448 16823 4450
rect 14365 4392 14370 4448
rect 14426 4392 16762 4448
rect 16818 4392 16823 4448
rect 14365 4390 16823 4392
rect 14365 4387 14431 4390
rect 16757 4387 16823 4390
rect 4825 4384 5141 4385
rect 4825 4320 4831 4384
rect 4895 4320 4911 4384
rect 4975 4320 4991 4384
rect 5055 4320 5071 4384
rect 5135 4320 5141 4384
rect 4825 4319 5141 4320
rect 11264 4384 11580 4385
rect 11264 4320 11270 4384
rect 11334 4320 11350 4384
rect 11414 4320 11430 4384
rect 11494 4320 11510 4384
rect 11574 4320 11580 4384
rect 11264 4319 11580 4320
rect 17703 4384 18019 4385
rect 17703 4320 17709 4384
rect 17773 4320 17789 4384
rect 17853 4320 17869 4384
rect 17933 4320 17949 4384
rect 18013 4320 18019 4384
rect 17703 4319 18019 4320
rect 24142 4384 24458 4385
rect 24142 4320 24148 4384
rect 24212 4320 24228 4384
rect 24292 4320 24308 4384
rect 24372 4320 24388 4384
rect 24452 4320 24458 4384
rect 24142 4319 24458 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 16113 4042 16179 4045
rect 17769 4042 17835 4045
rect 16113 4040 17835 4042
rect 16113 3984 16118 4040
rect 16174 3984 17774 4040
rect 17830 3984 17835 4040
rect 16113 3982 17835 3984
rect 16113 3979 16179 3982
rect 17769 3979 17835 3982
rect 26509 3906 26575 3909
rect 27188 3906 27988 3936
rect 26509 3904 27988 3906
rect 26509 3848 26514 3904
rect 26570 3848 27988 3904
rect 26509 3846 27988 3848
rect 26509 3843 26575 3846
rect 4165 3840 4481 3841
rect 4165 3776 4171 3840
rect 4235 3776 4251 3840
rect 4315 3776 4331 3840
rect 4395 3776 4411 3840
rect 4475 3776 4481 3840
rect 4165 3775 4481 3776
rect 10604 3840 10920 3841
rect 10604 3776 10610 3840
rect 10674 3776 10690 3840
rect 10754 3776 10770 3840
rect 10834 3776 10850 3840
rect 10914 3776 10920 3840
rect 10604 3775 10920 3776
rect 17043 3840 17359 3841
rect 17043 3776 17049 3840
rect 17113 3776 17129 3840
rect 17193 3776 17209 3840
rect 17273 3776 17289 3840
rect 17353 3776 17359 3840
rect 17043 3775 17359 3776
rect 23482 3840 23798 3841
rect 23482 3776 23488 3840
rect 23552 3776 23568 3840
rect 23632 3776 23648 3840
rect 23712 3776 23728 3840
rect 23792 3776 23798 3840
rect 27188 3816 27988 3846
rect 23482 3775 23798 3776
rect 4825 3296 5141 3297
rect 4825 3232 4831 3296
rect 4895 3232 4911 3296
rect 4975 3232 4991 3296
rect 5055 3232 5071 3296
rect 5135 3232 5141 3296
rect 4825 3231 5141 3232
rect 11264 3296 11580 3297
rect 11264 3232 11270 3296
rect 11334 3232 11350 3296
rect 11414 3232 11430 3296
rect 11494 3232 11510 3296
rect 11574 3232 11580 3296
rect 11264 3231 11580 3232
rect 17703 3296 18019 3297
rect 17703 3232 17709 3296
rect 17773 3232 17789 3296
rect 17853 3232 17869 3296
rect 17933 3232 17949 3296
rect 18013 3232 18019 3296
rect 17703 3231 18019 3232
rect 24142 3296 24458 3297
rect 24142 3232 24148 3296
rect 24212 3232 24228 3296
rect 24292 3232 24308 3296
rect 24372 3232 24388 3296
rect 24452 3232 24458 3296
rect 24142 3231 24458 3232
rect 4165 2752 4481 2753
rect 4165 2688 4171 2752
rect 4235 2688 4251 2752
rect 4315 2688 4331 2752
rect 4395 2688 4411 2752
rect 4475 2688 4481 2752
rect 4165 2687 4481 2688
rect 10604 2752 10920 2753
rect 10604 2688 10610 2752
rect 10674 2688 10690 2752
rect 10754 2688 10770 2752
rect 10834 2688 10850 2752
rect 10914 2688 10920 2752
rect 10604 2687 10920 2688
rect 17043 2752 17359 2753
rect 17043 2688 17049 2752
rect 17113 2688 17129 2752
rect 17193 2688 17209 2752
rect 17273 2688 17289 2752
rect 17353 2688 17359 2752
rect 17043 2687 17359 2688
rect 23482 2752 23798 2753
rect 23482 2688 23488 2752
rect 23552 2688 23568 2752
rect 23632 2688 23648 2752
rect 23712 2688 23728 2752
rect 23792 2688 23798 2752
rect 23482 2687 23798 2688
rect 4825 2208 5141 2209
rect 4825 2144 4831 2208
rect 4895 2144 4911 2208
rect 4975 2144 4991 2208
rect 5055 2144 5071 2208
rect 5135 2144 5141 2208
rect 4825 2143 5141 2144
rect 11264 2208 11580 2209
rect 11264 2144 11270 2208
rect 11334 2144 11350 2208
rect 11414 2144 11430 2208
rect 11494 2144 11510 2208
rect 11574 2144 11580 2208
rect 11264 2143 11580 2144
rect 17703 2208 18019 2209
rect 17703 2144 17709 2208
rect 17773 2144 17789 2208
rect 17853 2144 17869 2208
rect 17933 2144 17949 2208
rect 18013 2144 18019 2208
rect 17703 2143 18019 2144
rect 24142 2208 24458 2209
rect 24142 2144 24148 2208
rect 24212 2144 24228 2208
rect 24292 2144 24308 2208
rect 24372 2144 24388 2208
rect 24452 2144 24458 2208
rect 24142 2143 24458 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
<< via3 >>
rect 4171 27772 4235 27776
rect 4171 27716 4175 27772
rect 4175 27716 4231 27772
rect 4231 27716 4235 27772
rect 4171 27712 4235 27716
rect 4251 27772 4315 27776
rect 4251 27716 4255 27772
rect 4255 27716 4311 27772
rect 4311 27716 4315 27772
rect 4251 27712 4315 27716
rect 4331 27772 4395 27776
rect 4331 27716 4335 27772
rect 4335 27716 4391 27772
rect 4391 27716 4395 27772
rect 4331 27712 4395 27716
rect 4411 27772 4475 27776
rect 4411 27716 4415 27772
rect 4415 27716 4471 27772
rect 4471 27716 4475 27772
rect 4411 27712 4475 27716
rect 10610 27772 10674 27776
rect 10610 27716 10614 27772
rect 10614 27716 10670 27772
rect 10670 27716 10674 27772
rect 10610 27712 10674 27716
rect 10690 27772 10754 27776
rect 10690 27716 10694 27772
rect 10694 27716 10750 27772
rect 10750 27716 10754 27772
rect 10690 27712 10754 27716
rect 10770 27772 10834 27776
rect 10770 27716 10774 27772
rect 10774 27716 10830 27772
rect 10830 27716 10834 27772
rect 10770 27712 10834 27716
rect 10850 27772 10914 27776
rect 10850 27716 10854 27772
rect 10854 27716 10910 27772
rect 10910 27716 10914 27772
rect 10850 27712 10914 27716
rect 17049 27772 17113 27776
rect 17049 27716 17053 27772
rect 17053 27716 17109 27772
rect 17109 27716 17113 27772
rect 17049 27712 17113 27716
rect 17129 27772 17193 27776
rect 17129 27716 17133 27772
rect 17133 27716 17189 27772
rect 17189 27716 17193 27772
rect 17129 27712 17193 27716
rect 17209 27772 17273 27776
rect 17209 27716 17213 27772
rect 17213 27716 17269 27772
rect 17269 27716 17273 27772
rect 17209 27712 17273 27716
rect 17289 27772 17353 27776
rect 17289 27716 17293 27772
rect 17293 27716 17349 27772
rect 17349 27716 17353 27772
rect 17289 27712 17353 27716
rect 23488 27772 23552 27776
rect 23488 27716 23492 27772
rect 23492 27716 23548 27772
rect 23548 27716 23552 27772
rect 23488 27712 23552 27716
rect 23568 27772 23632 27776
rect 23568 27716 23572 27772
rect 23572 27716 23628 27772
rect 23628 27716 23632 27772
rect 23568 27712 23632 27716
rect 23648 27772 23712 27776
rect 23648 27716 23652 27772
rect 23652 27716 23708 27772
rect 23708 27716 23712 27772
rect 23648 27712 23712 27716
rect 23728 27772 23792 27776
rect 23728 27716 23732 27772
rect 23732 27716 23788 27772
rect 23788 27716 23792 27772
rect 23728 27712 23792 27716
rect 4831 27228 4895 27232
rect 4831 27172 4835 27228
rect 4835 27172 4891 27228
rect 4891 27172 4895 27228
rect 4831 27168 4895 27172
rect 4911 27228 4975 27232
rect 4911 27172 4915 27228
rect 4915 27172 4971 27228
rect 4971 27172 4975 27228
rect 4911 27168 4975 27172
rect 4991 27228 5055 27232
rect 4991 27172 4995 27228
rect 4995 27172 5051 27228
rect 5051 27172 5055 27228
rect 4991 27168 5055 27172
rect 5071 27228 5135 27232
rect 5071 27172 5075 27228
rect 5075 27172 5131 27228
rect 5131 27172 5135 27228
rect 5071 27168 5135 27172
rect 11270 27228 11334 27232
rect 11270 27172 11274 27228
rect 11274 27172 11330 27228
rect 11330 27172 11334 27228
rect 11270 27168 11334 27172
rect 11350 27228 11414 27232
rect 11350 27172 11354 27228
rect 11354 27172 11410 27228
rect 11410 27172 11414 27228
rect 11350 27168 11414 27172
rect 11430 27228 11494 27232
rect 11430 27172 11434 27228
rect 11434 27172 11490 27228
rect 11490 27172 11494 27228
rect 11430 27168 11494 27172
rect 11510 27228 11574 27232
rect 11510 27172 11514 27228
rect 11514 27172 11570 27228
rect 11570 27172 11574 27228
rect 11510 27168 11574 27172
rect 17709 27228 17773 27232
rect 17709 27172 17713 27228
rect 17713 27172 17769 27228
rect 17769 27172 17773 27228
rect 17709 27168 17773 27172
rect 17789 27228 17853 27232
rect 17789 27172 17793 27228
rect 17793 27172 17849 27228
rect 17849 27172 17853 27228
rect 17789 27168 17853 27172
rect 17869 27228 17933 27232
rect 17869 27172 17873 27228
rect 17873 27172 17929 27228
rect 17929 27172 17933 27228
rect 17869 27168 17933 27172
rect 17949 27228 18013 27232
rect 17949 27172 17953 27228
rect 17953 27172 18009 27228
rect 18009 27172 18013 27228
rect 17949 27168 18013 27172
rect 24148 27228 24212 27232
rect 24148 27172 24152 27228
rect 24152 27172 24208 27228
rect 24208 27172 24212 27228
rect 24148 27168 24212 27172
rect 24228 27228 24292 27232
rect 24228 27172 24232 27228
rect 24232 27172 24288 27228
rect 24288 27172 24292 27228
rect 24228 27168 24292 27172
rect 24308 27228 24372 27232
rect 24308 27172 24312 27228
rect 24312 27172 24368 27228
rect 24368 27172 24372 27228
rect 24308 27168 24372 27172
rect 24388 27228 24452 27232
rect 24388 27172 24392 27228
rect 24392 27172 24448 27228
rect 24448 27172 24452 27228
rect 24388 27168 24452 27172
rect 4171 26684 4235 26688
rect 4171 26628 4175 26684
rect 4175 26628 4231 26684
rect 4231 26628 4235 26684
rect 4171 26624 4235 26628
rect 4251 26684 4315 26688
rect 4251 26628 4255 26684
rect 4255 26628 4311 26684
rect 4311 26628 4315 26684
rect 4251 26624 4315 26628
rect 4331 26684 4395 26688
rect 4331 26628 4335 26684
rect 4335 26628 4391 26684
rect 4391 26628 4395 26684
rect 4331 26624 4395 26628
rect 4411 26684 4475 26688
rect 4411 26628 4415 26684
rect 4415 26628 4471 26684
rect 4471 26628 4475 26684
rect 4411 26624 4475 26628
rect 10610 26684 10674 26688
rect 10610 26628 10614 26684
rect 10614 26628 10670 26684
rect 10670 26628 10674 26684
rect 10610 26624 10674 26628
rect 10690 26684 10754 26688
rect 10690 26628 10694 26684
rect 10694 26628 10750 26684
rect 10750 26628 10754 26684
rect 10690 26624 10754 26628
rect 10770 26684 10834 26688
rect 10770 26628 10774 26684
rect 10774 26628 10830 26684
rect 10830 26628 10834 26684
rect 10770 26624 10834 26628
rect 10850 26684 10914 26688
rect 10850 26628 10854 26684
rect 10854 26628 10910 26684
rect 10910 26628 10914 26684
rect 10850 26624 10914 26628
rect 17049 26684 17113 26688
rect 17049 26628 17053 26684
rect 17053 26628 17109 26684
rect 17109 26628 17113 26684
rect 17049 26624 17113 26628
rect 17129 26684 17193 26688
rect 17129 26628 17133 26684
rect 17133 26628 17189 26684
rect 17189 26628 17193 26684
rect 17129 26624 17193 26628
rect 17209 26684 17273 26688
rect 17209 26628 17213 26684
rect 17213 26628 17269 26684
rect 17269 26628 17273 26684
rect 17209 26624 17273 26628
rect 17289 26684 17353 26688
rect 17289 26628 17293 26684
rect 17293 26628 17349 26684
rect 17349 26628 17353 26684
rect 17289 26624 17353 26628
rect 23488 26684 23552 26688
rect 23488 26628 23492 26684
rect 23492 26628 23548 26684
rect 23548 26628 23552 26684
rect 23488 26624 23552 26628
rect 23568 26684 23632 26688
rect 23568 26628 23572 26684
rect 23572 26628 23628 26684
rect 23628 26628 23632 26684
rect 23568 26624 23632 26628
rect 23648 26684 23712 26688
rect 23648 26628 23652 26684
rect 23652 26628 23708 26684
rect 23708 26628 23712 26684
rect 23648 26624 23712 26628
rect 23728 26684 23792 26688
rect 23728 26628 23732 26684
rect 23732 26628 23788 26684
rect 23788 26628 23792 26684
rect 23728 26624 23792 26628
rect 4831 26140 4895 26144
rect 4831 26084 4835 26140
rect 4835 26084 4891 26140
rect 4891 26084 4895 26140
rect 4831 26080 4895 26084
rect 4911 26140 4975 26144
rect 4911 26084 4915 26140
rect 4915 26084 4971 26140
rect 4971 26084 4975 26140
rect 4911 26080 4975 26084
rect 4991 26140 5055 26144
rect 4991 26084 4995 26140
rect 4995 26084 5051 26140
rect 5051 26084 5055 26140
rect 4991 26080 5055 26084
rect 5071 26140 5135 26144
rect 5071 26084 5075 26140
rect 5075 26084 5131 26140
rect 5131 26084 5135 26140
rect 5071 26080 5135 26084
rect 11270 26140 11334 26144
rect 11270 26084 11274 26140
rect 11274 26084 11330 26140
rect 11330 26084 11334 26140
rect 11270 26080 11334 26084
rect 11350 26140 11414 26144
rect 11350 26084 11354 26140
rect 11354 26084 11410 26140
rect 11410 26084 11414 26140
rect 11350 26080 11414 26084
rect 11430 26140 11494 26144
rect 11430 26084 11434 26140
rect 11434 26084 11490 26140
rect 11490 26084 11494 26140
rect 11430 26080 11494 26084
rect 11510 26140 11574 26144
rect 11510 26084 11514 26140
rect 11514 26084 11570 26140
rect 11570 26084 11574 26140
rect 11510 26080 11574 26084
rect 17709 26140 17773 26144
rect 17709 26084 17713 26140
rect 17713 26084 17769 26140
rect 17769 26084 17773 26140
rect 17709 26080 17773 26084
rect 17789 26140 17853 26144
rect 17789 26084 17793 26140
rect 17793 26084 17849 26140
rect 17849 26084 17853 26140
rect 17789 26080 17853 26084
rect 17869 26140 17933 26144
rect 17869 26084 17873 26140
rect 17873 26084 17929 26140
rect 17929 26084 17933 26140
rect 17869 26080 17933 26084
rect 17949 26140 18013 26144
rect 17949 26084 17953 26140
rect 17953 26084 18009 26140
rect 18009 26084 18013 26140
rect 17949 26080 18013 26084
rect 24148 26140 24212 26144
rect 24148 26084 24152 26140
rect 24152 26084 24208 26140
rect 24208 26084 24212 26140
rect 24148 26080 24212 26084
rect 24228 26140 24292 26144
rect 24228 26084 24232 26140
rect 24232 26084 24288 26140
rect 24288 26084 24292 26140
rect 24228 26080 24292 26084
rect 24308 26140 24372 26144
rect 24308 26084 24312 26140
rect 24312 26084 24368 26140
rect 24368 26084 24372 26140
rect 24308 26080 24372 26084
rect 24388 26140 24452 26144
rect 24388 26084 24392 26140
rect 24392 26084 24448 26140
rect 24448 26084 24452 26140
rect 24388 26080 24452 26084
rect 4171 25596 4235 25600
rect 4171 25540 4175 25596
rect 4175 25540 4231 25596
rect 4231 25540 4235 25596
rect 4171 25536 4235 25540
rect 4251 25596 4315 25600
rect 4251 25540 4255 25596
rect 4255 25540 4311 25596
rect 4311 25540 4315 25596
rect 4251 25536 4315 25540
rect 4331 25596 4395 25600
rect 4331 25540 4335 25596
rect 4335 25540 4391 25596
rect 4391 25540 4395 25596
rect 4331 25536 4395 25540
rect 4411 25596 4475 25600
rect 4411 25540 4415 25596
rect 4415 25540 4471 25596
rect 4471 25540 4475 25596
rect 4411 25536 4475 25540
rect 10610 25596 10674 25600
rect 10610 25540 10614 25596
rect 10614 25540 10670 25596
rect 10670 25540 10674 25596
rect 10610 25536 10674 25540
rect 10690 25596 10754 25600
rect 10690 25540 10694 25596
rect 10694 25540 10750 25596
rect 10750 25540 10754 25596
rect 10690 25536 10754 25540
rect 10770 25596 10834 25600
rect 10770 25540 10774 25596
rect 10774 25540 10830 25596
rect 10830 25540 10834 25596
rect 10770 25536 10834 25540
rect 10850 25596 10914 25600
rect 10850 25540 10854 25596
rect 10854 25540 10910 25596
rect 10910 25540 10914 25596
rect 10850 25536 10914 25540
rect 17049 25596 17113 25600
rect 17049 25540 17053 25596
rect 17053 25540 17109 25596
rect 17109 25540 17113 25596
rect 17049 25536 17113 25540
rect 17129 25596 17193 25600
rect 17129 25540 17133 25596
rect 17133 25540 17189 25596
rect 17189 25540 17193 25596
rect 17129 25536 17193 25540
rect 17209 25596 17273 25600
rect 17209 25540 17213 25596
rect 17213 25540 17269 25596
rect 17269 25540 17273 25596
rect 17209 25536 17273 25540
rect 17289 25596 17353 25600
rect 17289 25540 17293 25596
rect 17293 25540 17349 25596
rect 17349 25540 17353 25596
rect 17289 25536 17353 25540
rect 23488 25596 23552 25600
rect 23488 25540 23492 25596
rect 23492 25540 23548 25596
rect 23548 25540 23552 25596
rect 23488 25536 23552 25540
rect 23568 25596 23632 25600
rect 23568 25540 23572 25596
rect 23572 25540 23628 25596
rect 23628 25540 23632 25596
rect 23568 25536 23632 25540
rect 23648 25596 23712 25600
rect 23648 25540 23652 25596
rect 23652 25540 23708 25596
rect 23708 25540 23712 25596
rect 23648 25536 23712 25540
rect 23728 25596 23792 25600
rect 23728 25540 23732 25596
rect 23732 25540 23788 25596
rect 23788 25540 23792 25596
rect 23728 25536 23792 25540
rect 4831 25052 4895 25056
rect 4831 24996 4835 25052
rect 4835 24996 4891 25052
rect 4891 24996 4895 25052
rect 4831 24992 4895 24996
rect 4911 25052 4975 25056
rect 4911 24996 4915 25052
rect 4915 24996 4971 25052
rect 4971 24996 4975 25052
rect 4911 24992 4975 24996
rect 4991 25052 5055 25056
rect 4991 24996 4995 25052
rect 4995 24996 5051 25052
rect 5051 24996 5055 25052
rect 4991 24992 5055 24996
rect 5071 25052 5135 25056
rect 5071 24996 5075 25052
rect 5075 24996 5131 25052
rect 5131 24996 5135 25052
rect 5071 24992 5135 24996
rect 11270 25052 11334 25056
rect 11270 24996 11274 25052
rect 11274 24996 11330 25052
rect 11330 24996 11334 25052
rect 11270 24992 11334 24996
rect 11350 25052 11414 25056
rect 11350 24996 11354 25052
rect 11354 24996 11410 25052
rect 11410 24996 11414 25052
rect 11350 24992 11414 24996
rect 11430 25052 11494 25056
rect 11430 24996 11434 25052
rect 11434 24996 11490 25052
rect 11490 24996 11494 25052
rect 11430 24992 11494 24996
rect 11510 25052 11574 25056
rect 11510 24996 11514 25052
rect 11514 24996 11570 25052
rect 11570 24996 11574 25052
rect 11510 24992 11574 24996
rect 17709 25052 17773 25056
rect 17709 24996 17713 25052
rect 17713 24996 17769 25052
rect 17769 24996 17773 25052
rect 17709 24992 17773 24996
rect 17789 25052 17853 25056
rect 17789 24996 17793 25052
rect 17793 24996 17849 25052
rect 17849 24996 17853 25052
rect 17789 24992 17853 24996
rect 17869 25052 17933 25056
rect 17869 24996 17873 25052
rect 17873 24996 17929 25052
rect 17929 24996 17933 25052
rect 17869 24992 17933 24996
rect 17949 25052 18013 25056
rect 17949 24996 17953 25052
rect 17953 24996 18009 25052
rect 18009 24996 18013 25052
rect 17949 24992 18013 24996
rect 24148 25052 24212 25056
rect 24148 24996 24152 25052
rect 24152 24996 24208 25052
rect 24208 24996 24212 25052
rect 24148 24992 24212 24996
rect 24228 25052 24292 25056
rect 24228 24996 24232 25052
rect 24232 24996 24288 25052
rect 24288 24996 24292 25052
rect 24228 24992 24292 24996
rect 24308 25052 24372 25056
rect 24308 24996 24312 25052
rect 24312 24996 24368 25052
rect 24368 24996 24372 25052
rect 24308 24992 24372 24996
rect 24388 25052 24452 25056
rect 24388 24996 24392 25052
rect 24392 24996 24448 25052
rect 24448 24996 24452 25052
rect 24388 24992 24452 24996
rect 4171 24508 4235 24512
rect 4171 24452 4175 24508
rect 4175 24452 4231 24508
rect 4231 24452 4235 24508
rect 4171 24448 4235 24452
rect 4251 24508 4315 24512
rect 4251 24452 4255 24508
rect 4255 24452 4311 24508
rect 4311 24452 4315 24508
rect 4251 24448 4315 24452
rect 4331 24508 4395 24512
rect 4331 24452 4335 24508
rect 4335 24452 4391 24508
rect 4391 24452 4395 24508
rect 4331 24448 4395 24452
rect 4411 24508 4475 24512
rect 4411 24452 4415 24508
rect 4415 24452 4471 24508
rect 4471 24452 4475 24508
rect 4411 24448 4475 24452
rect 10610 24508 10674 24512
rect 10610 24452 10614 24508
rect 10614 24452 10670 24508
rect 10670 24452 10674 24508
rect 10610 24448 10674 24452
rect 10690 24508 10754 24512
rect 10690 24452 10694 24508
rect 10694 24452 10750 24508
rect 10750 24452 10754 24508
rect 10690 24448 10754 24452
rect 10770 24508 10834 24512
rect 10770 24452 10774 24508
rect 10774 24452 10830 24508
rect 10830 24452 10834 24508
rect 10770 24448 10834 24452
rect 10850 24508 10914 24512
rect 10850 24452 10854 24508
rect 10854 24452 10910 24508
rect 10910 24452 10914 24508
rect 10850 24448 10914 24452
rect 17049 24508 17113 24512
rect 17049 24452 17053 24508
rect 17053 24452 17109 24508
rect 17109 24452 17113 24508
rect 17049 24448 17113 24452
rect 17129 24508 17193 24512
rect 17129 24452 17133 24508
rect 17133 24452 17189 24508
rect 17189 24452 17193 24508
rect 17129 24448 17193 24452
rect 17209 24508 17273 24512
rect 17209 24452 17213 24508
rect 17213 24452 17269 24508
rect 17269 24452 17273 24508
rect 17209 24448 17273 24452
rect 17289 24508 17353 24512
rect 17289 24452 17293 24508
rect 17293 24452 17349 24508
rect 17349 24452 17353 24508
rect 17289 24448 17353 24452
rect 23488 24508 23552 24512
rect 23488 24452 23492 24508
rect 23492 24452 23548 24508
rect 23548 24452 23552 24508
rect 23488 24448 23552 24452
rect 23568 24508 23632 24512
rect 23568 24452 23572 24508
rect 23572 24452 23628 24508
rect 23628 24452 23632 24508
rect 23568 24448 23632 24452
rect 23648 24508 23712 24512
rect 23648 24452 23652 24508
rect 23652 24452 23708 24508
rect 23708 24452 23712 24508
rect 23648 24448 23712 24452
rect 23728 24508 23792 24512
rect 23728 24452 23732 24508
rect 23732 24452 23788 24508
rect 23788 24452 23792 24508
rect 23728 24448 23792 24452
rect 4831 23964 4895 23968
rect 4831 23908 4835 23964
rect 4835 23908 4891 23964
rect 4891 23908 4895 23964
rect 4831 23904 4895 23908
rect 4911 23964 4975 23968
rect 4911 23908 4915 23964
rect 4915 23908 4971 23964
rect 4971 23908 4975 23964
rect 4911 23904 4975 23908
rect 4991 23964 5055 23968
rect 4991 23908 4995 23964
rect 4995 23908 5051 23964
rect 5051 23908 5055 23964
rect 4991 23904 5055 23908
rect 5071 23964 5135 23968
rect 5071 23908 5075 23964
rect 5075 23908 5131 23964
rect 5131 23908 5135 23964
rect 5071 23904 5135 23908
rect 11270 23964 11334 23968
rect 11270 23908 11274 23964
rect 11274 23908 11330 23964
rect 11330 23908 11334 23964
rect 11270 23904 11334 23908
rect 11350 23964 11414 23968
rect 11350 23908 11354 23964
rect 11354 23908 11410 23964
rect 11410 23908 11414 23964
rect 11350 23904 11414 23908
rect 11430 23964 11494 23968
rect 11430 23908 11434 23964
rect 11434 23908 11490 23964
rect 11490 23908 11494 23964
rect 11430 23904 11494 23908
rect 11510 23964 11574 23968
rect 11510 23908 11514 23964
rect 11514 23908 11570 23964
rect 11570 23908 11574 23964
rect 11510 23904 11574 23908
rect 17709 23964 17773 23968
rect 17709 23908 17713 23964
rect 17713 23908 17769 23964
rect 17769 23908 17773 23964
rect 17709 23904 17773 23908
rect 17789 23964 17853 23968
rect 17789 23908 17793 23964
rect 17793 23908 17849 23964
rect 17849 23908 17853 23964
rect 17789 23904 17853 23908
rect 17869 23964 17933 23968
rect 17869 23908 17873 23964
rect 17873 23908 17929 23964
rect 17929 23908 17933 23964
rect 17869 23904 17933 23908
rect 17949 23964 18013 23968
rect 17949 23908 17953 23964
rect 17953 23908 18009 23964
rect 18009 23908 18013 23964
rect 17949 23904 18013 23908
rect 24148 23964 24212 23968
rect 24148 23908 24152 23964
rect 24152 23908 24208 23964
rect 24208 23908 24212 23964
rect 24148 23904 24212 23908
rect 24228 23964 24292 23968
rect 24228 23908 24232 23964
rect 24232 23908 24288 23964
rect 24288 23908 24292 23964
rect 24228 23904 24292 23908
rect 24308 23964 24372 23968
rect 24308 23908 24312 23964
rect 24312 23908 24368 23964
rect 24368 23908 24372 23964
rect 24308 23904 24372 23908
rect 24388 23964 24452 23968
rect 24388 23908 24392 23964
rect 24392 23908 24448 23964
rect 24448 23908 24452 23964
rect 24388 23904 24452 23908
rect 4171 23420 4235 23424
rect 4171 23364 4175 23420
rect 4175 23364 4231 23420
rect 4231 23364 4235 23420
rect 4171 23360 4235 23364
rect 4251 23420 4315 23424
rect 4251 23364 4255 23420
rect 4255 23364 4311 23420
rect 4311 23364 4315 23420
rect 4251 23360 4315 23364
rect 4331 23420 4395 23424
rect 4331 23364 4335 23420
rect 4335 23364 4391 23420
rect 4391 23364 4395 23420
rect 4331 23360 4395 23364
rect 4411 23420 4475 23424
rect 4411 23364 4415 23420
rect 4415 23364 4471 23420
rect 4471 23364 4475 23420
rect 4411 23360 4475 23364
rect 10610 23420 10674 23424
rect 10610 23364 10614 23420
rect 10614 23364 10670 23420
rect 10670 23364 10674 23420
rect 10610 23360 10674 23364
rect 10690 23420 10754 23424
rect 10690 23364 10694 23420
rect 10694 23364 10750 23420
rect 10750 23364 10754 23420
rect 10690 23360 10754 23364
rect 10770 23420 10834 23424
rect 10770 23364 10774 23420
rect 10774 23364 10830 23420
rect 10830 23364 10834 23420
rect 10770 23360 10834 23364
rect 10850 23420 10914 23424
rect 10850 23364 10854 23420
rect 10854 23364 10910 23420
rect 10910 23364 10914 23420
rect 10850 23360 10914 23364
rect 17049 23420 17113 23424
rect 17049 23364 17053 23420
rect 17053 23364 17109 23420
rect 17109 23364 17113 23420
rect 17049 23360 17113 23364
rect 17129 23420 17193 23424
rect 17129 23364 17133 23420
rect 17133 23364 17189 23420
rect 17189 23364 17193 23420
rect 17129 23360 17193 23364
rect 17209 23420 17273 23424
rect 17209 23364 17213 23420
rect 17213 23364 17269 23420
rect 17269 23364 17273 23420
rect 17209 23360 17273 23364
rect 17289 23420 17353 23424
rect 17289 23364 17293 23420
rect 17293 23364 17349 23420
rect 17349 23364 17353 23420
rect 17289 23360 17353 23364
rect 23488 23420 23552 23424
rect 23488 23364 23492 23420
rect 23492 23364 23548 23420
rect 23548 23364 23552 23420
rect 23488 23360 23552 23364
rect 23568 23420 23632 23424
rect 23568 23364 23572 23420
rect 23572 23364 23628 23420
rect 23628 23364 23632 23420
rect 23568 23360 23632 23364
rect 23648 23420 23712 23424
rect 23648 23364 23652 23420
rect 23652 23364 23708 23420
rect 23708 23364 23712 23420
rect 23648 23360 23712 23364
rect 23728 23420 23792 23424
rect 23728 23364 23732 23420
rect 23732 23364 23788 23420
rect 23788 23364 23792 23420
rect 23728 23360 23792 23364
rect 4831 22876 4895 22880
rect 4831 22820 4835 22876
rect 4835 22820 4891 22876
rect 4891 22820 4895 22876
rect 4831 22816 4895 22820
rect 4911 22876 4975 22880
rect 4911 22820 4915 22876
rect 4915 22820 4971 22876
rect 4971 22820 4975 22876
rect 4911 22816 4975 22820
rect 4991 22876 5055 22880
rect 4991 22820 4995 22876
rect 4995 22820 5051 22876
rect 5051 22820 5055 22876
rect 4991 22816 5055 22820
rect 5071 22876 5135 22880
rect 5071 22820 5075 22876
rect 5075 22820 5131 22876
rect 5131 22820 5135 22876
rect 5071 22816 5135 22820
rect 11270 22876 11334 22880
rect 11270 22820 11274 22876
rect 11274 22820 11330 22876
rect 11330 22820 11334 22876
rect 11270 22816 11334 22820
rect 11350 22876 11414 22880
rect 11350 22820 11354 22876
rect 11354 22820 11410 22876
rect 11410 22820 11414 22876
rect 11350 22816 11414 22820
rect 11430 22876 11494 22880
rect 11430 22820 11434 22876
rect 11434 22820 11490 22876
rect 11490 22820 11494 22876
rect 11430 22816 11494 22820
rect 11510 22876 11574 22880
rect 11510 22820 11514 22876
rect 11514 22820 11570 22876
rect 11570 22820 11574 22876
rect 11510 22816 11574 22820
rect 17709 22876 17773 22880
rect 17709 22820 17713 22876
rect 17713 22820 17769 22876
rect 17769 22820 17773 22876
rect 17709 22816 17773 22820
rect 17789 22876 17853 22880
rect 17789 22820 17793 22876
rect 17793 22820 17849 22876
rect 17849 22820 17853 22876
rect 17789 22816 17853 22820
rect 17869 22876 17933 22880
rect 17869 22820 17873 22876
rect 17873 22820 17929 22876
rect 17929 22820 17933 22876
rect 17869 22816 17933 22820
rect 17949 22876 18013 22880
rect 17949 22820 17953 22876
rect 17953 22820 18009 22876
rect 18009 22820 18013 22876
rect 17949 22816 18013 22820
rect 24148 22876 24212 22880
rect 24148 22820 24152 22876
rect 24152 22820 24208 22876
rect 24208 22820 24212 22876
rect 24148 22816 24212 22820
rect 24228 22876 24292 22880
rect 24228 22820 24232 22876
rect 24232 22820 24288 22876
rect 24288 22820 24292 22876
rect 24228 22816 24292 22820
rect 24308 22876 24372 22880
rect 24308 22820 24312 22876
rect 24312 22820 24368 22876
rect 24368 22820 24372 22876
rect 24308 22816 24372 22820
rect 24388 22876 24452 22880
rect 24388 22820 24392 22876
rect 24392 22820 24448 22876
rect 24448 22820 24452 22876
rect 24388 22816 24452 22820
rect 4171 22332 4235 22336
rect 4171 22276 4175 22332
rect 4175 22276 4231 22332
rect 4231 22276 4235 22332
rect 4171 22272 4235 22276
rect 4251 22332 4315 22336
rect 4251 22276 4255 22332
rect 4255 22276 4311 22332
rect 4311 22276 4315 22332
rect 4251 22272 4315 22276
rect 4331 22332 4395 22336
rect 4331 22276 4335 22332
rect 4335 22276 4391 22332
rect 4391 22276 4395 22332
rect 4331 22272 4395 22276
rect 4411 22332 4475 22336
rect 4411 22276 4415 22332
rect 4415 22276 4471 22332
rect 4471 22276 4475 22332
rect 4411 22272 4475 22276
rect 10610 22332 10674 22336
rect 10610 22276 10614 22332
rect 10614 22276 10670 22332
rect 10670 22276 10674 22332
rect 10610 22272 10674 22276
rect 10690 22332 10754 22336
rect 10690 22276 10694 22332
rect 10694 22276 10750 22332
rect 10750 22276 10754 22332
rect 10690 22272 10754 22276
rect 10770 22332 10834 22336
rect 10770 22276 10774 22332
rect 10774 22276 10830 22332
rect 10830 22276 10834 22332
rect 10770 22272 10834 22276
rect 10850 22332 10914 22336
rect 10850 22276 10854 22332
rect 10854 22276 10910 22332
rect 10910 22276 10914 22332
rect 10850 22272 10914 22276
rect 17049 22332 17113 22336
rect 17049 22276 17053 22332
rect 17053 22276 17109 22332
rect 17109 22276 17113 22332
rect 17049 22272 17113 22276
rect 17129 22332 17193 22336
rect 17129 22276 17133 22332
rect 17133 22276 17189 22332
rect 17189 22276 17193 22332
rect 17129 22272 17193 22276
rect 17209 22332 17273 22336
rect 17209 22276 17213 22332
rect 17213 22276 17269 22332
rect 17269 22276 17273 22332
rect 17209 22272 17273 22276
rect 17289 22332 17353 22336
rect 17289 22276 17293 22332
rect 17293 22276 17349 22332
rect 17349 22276 17353 22332
rect 17289 22272 17353 22276
rect 23488 22332 23552 22336
rect 23488 22276 23492 22332
rect 23492 22276 23548 22332
rect 23548 22276 23552 22332
rect 23488 22272 23552 22276
rect 23568 22332 23632 22336
rect 23568 22276 23572 22332
rect 23572 22276 23628 22332
rect 23628 22276 23632 22332
rect 23568 22272 23632 22276
rect 23648 22332 23712 22336
rect 23648 22276 23652 22332
rect 23652 22276 23708 22332
rect 23708 22276 23712 22332
rect 23648 22272 23712 22276
rect 23728 22332 23792 22336
rect 23728 22276 23732 22332
rect 23732 22276 23788 22332
rect 23788 22276 23792 22332
rect 23728 22272 23792 22276
rect 4831 21788 4895 21792
rect 4831 21732 4835 21788
rect 4835 21732 4891 21788
rect 4891 21732 4895 21788
rect 4831 21728 4895 21732
rect 4911 21788 4975 21792
rect 4911 21732 4915 21788
rect 4915 21732 4971 21788
rect 4971 21732 4975 21788
rect 4911 21728 4975 21732
rect 4991 21788 5055 21792
rect 4991 21732 4995 21788
rect 4995 21732 5051 21788
rect 5051 21732 5055 21788
rect 4991 21728 5055 21732
rect 5071 21788 5135 21792
rect 5071 21732 5075 21788
rect 5075 21732 5131 21788
rect 5131 21732 5135 21788
rect 5071 21728 5135 21732
rect 11270 21788 11334 21792
rect 11270 21732 11274 21788
rect 11274 21732 11330 21788
rect 11330 21732 11334 21788
rect 11270 21728 11334 21732
rect 11350 21788 11414 21792
rect 11350 21732 11354 21788
rect 11354 21732 11410 21788
rect 11410 21732 11414 21788
rect 11350 21728 11414 21732
rect 11430 21788 11494 21792
rect 11430 21732 11434 21788
rect 11434 21732 11490 21788
rect 11490 21732 11494 21788
rect 11430 21728 11494 21732
rect 11510 21788 11574 21792
rect 11510 21732 11514 21788
rect 11514 21732 11570 21788
rect 11570 21732 11574 21788
rect 11510 21728 11574 21732
rect 17709 21788 17773 21792
rect 17709 21732 17713 21788
rect 17713 21732 17769 21788
rect 17769 21732 17773 21788
rect 17709 21728 17773 21732
rect 17789 21788 17853 21792
rect 17789 21732 17793 21788
rect 17793 21732 17849 21788
rect 17849 21732 17853 21788
rect 17789 21728 17853 21732
rect 17869 21788 17933 21792
rect 17869 21732 17873 21788
rect 17873 21732 17929 21788
rect 17929 21732 17933 21788
rect 17869 21728 17933 21732
rect 17949 21788 18013 21792
rect 17949 21732 17953 21788
rect 17953 21732 18009 21788
rect 18009 21732 18013 21788
rect 17949 21728 18013 21732
rect 24148 21788 24212 21792
rect 24148 21732 24152 21788
rect 24152 21732 24208 21788
rect 24208 21732 24212 21788
rect 24148 21728 24212 21732
rect 24228 21788 24292 21792
rect 24228 21732 24232 21788
rect 24232 21732 24288 21788
rect 24288 21732 24292 21788
rect 24228 21728 24292 21732
rect 24308 21788 24372 21792
rect 24308 21732 24312 21788
rect 24312 21732 24368 21788
rect 24368 21732 24372 21788
rect 24308 21728 24372 21732
rect 24388 21788 24452 21792
rect 24388 21732 24392 21788
rect 24392 21732 24448 21788
rect 24448 21732 24452 21788
rect 24388 21728 24452 21732
rect 4171 21244 4235 21248
rect 4171 21188 4175 21244
rect 4175 21188 4231 21244
rect 4231 21188 4235 21244
rect 4171 21184 4235 21188
rect 4251 21244 4315 21248
rect 4251 21188 4255 21244
rect 4255 21188 4311 21244
rect 4311 21188 4315 21244
rect 4251 21184 4315 21188
rect 4331 21244 4395 21248
rect 4331 21188 4335 21244
rect 4335 21188 4391 21244
rect 4391 21188 4395 21244
rect 4331 21184 4395 21188
rect 4411 21244 4475 21248
rect 4411 21188 4415 21244
rect 4415 21188 4471 21244
rect 4471 21188 4475 21244
rect 4411 21184 4475 21188
rect 10610 21244 10674 21248
rect 10610 21188 10614 21244
rect 10614 21188 10670 21244
rect 10670 21188 10674 21244
rect 10610 21184 10674 21188
rect 10690 21244 10754 21248
rect 10690 21188 10694 21244
rect 10694 21188 10750 21244
rect 10750 21188 10754 21244
rect 10690 21184 10754 21188
rect 10770 21244 10834 21248
rect 10770 21188 10774 21244
rect 10774 21188 10830 21244
rect 10830 21188 10834 21244
rect 10770 21184 10834 21188
rect 10850 21244 10914 21248
rect 10850 21188 10854 21244
rect 10854 21188 10910 21244
rect 10910 21188 10914 21244
rect 10850 21184 10914 21188
rect 17049 21244 17113 21248
rect 17049 21188 17053 21244
rect 17053 21188 17109 21244
rect 17109 21188 17113 21244
rect 17049 21184 17113 21188
rect 17129 21244 17193 21248
rect 17129 21188 17133 21244
rect 17133 21188 17189 21244
rect 17189 21188 17193 21244
rect 17129 21184 17193 21188
rect 17209 21244 17273 21248
rect 17209 21188 17213 21244
rect 17213 21188 17269 21244
rect 17269 21188 17273 21244
rect 17209 21184 17273 21188
rect 17289 21244 17353 21248
rect 17289 21188 17293 21244
rect 17293 21188 17349 21244
rect 17349 21188 17353 21244
rect 17289 21184 17353 21188
rect 23488 21244 23552 21248
rect 23488 21188 23492 21244
rect 23492 21188 23548 21244
rect 23548 21188 23552 21244
rect 23488 21184 23552 21188
rect 23568 21244 23632 21248
rect 23568 21188 23572 21244
rect 23572 21188 23628 21244
rect 23628 21188 23632 21244
rect 23568 21184 23632 21188
rect 23648 21244 23712 21248
rect 23648 21188 23652 21244
rect 23652 21188 23708 21244
rect 23708 21188 23712 21244
rect 23648 21184 23712 21188
rect 23728 21244 23792 21248
rect 23728 21188 23732 21244
rect 23732 21188 23788 21244
rect 23788 21188 23792 21244
rect 23728 21184 23792 21188
rect 15332 20708 15396 20772
rect 4831 20700 4895 20704
rect 4831 20644 4835 20700
rect 4835 20644 4891 20700
rect 4891 20644 4895 20700
rect 4831 20640 4895 20644
rect 4911 20700 4975 20704
rect 4911 20644 4915 20700
rect 4915 20644 4971 20700
rect 4971 20644 4975 20700
rect 4911 20640 4975 20644
rect 4991 20700 5055 20704
rect 4991 20644 4995 20700
rect 4995 20644 5051 20700
rect 5051 20644 5055 20700
rect 4991 20640 5055 20644
rect 5071 20700 5135 20704
rect 5071 20644 5075 20700
rect 5075 20644 5131 20700
rect 5131 20644 5135 20700
rect 5071 20640 5135 20644
rect 11270 20700 11334 20704
rect 11270 20644 11274 20700
rect 11274 20644 11330 20700
rect 11330 20644 11334 20700
rect 11270 20640 11334 20644
rect 11350 20700 11414 20704
rect 11350 20644 11354 20700
rect 11354 20644 11410 20700
rect 11410 20644 11414 20700
rect 11350 20640 11414 20644
rect 11430 20700 11494 20704
rect 11430 20644 11434 20700
rect 11434 20644 11490 20700
rect 11490 20644 11494 20700
rect 11430 20640 11494 20644
rect 11510 20700 11574 20704
rect 11510 20644 11514 20700
rect 11514 20644 11570 20700
rect 11570 20644 11574 20700
rect 11510 20640 11574 20644
rect 17709 20700 17773 20704
rect 17709 20644 17713 20700
rect 17713 20644 17769 20700
rect 17769 20644 17773 20700
rect 17709 20640 17773 20644
rect 17789 20700 17853 20704
rect 17789 20644 17793 20700
rect 17793 20644 17849 20700
rect 17849 20644 17853 20700
rect 17789 20640 17853 20644
rect 17869 20700 17933 20704
rect 17869 20644 17873 20700
rect 17873 20644 17929 20700
rect 17929 20644 17933 20700
rect 17869 20640 17933 20644
rect 17949 20700 18013 20704
rect 17949 20644 17953 20700
rect 17953 20644 18009 20700
rect 18009 20644 18013 20700
rect 17949 20640 18013 20644
rect 24148 20700 24212 20704
rect 24148 20644 24152 20700
rect 24152 20644 24208 20700
rect 24208 20644 24212 20700
rect 24148 20640 24212 20644
rect 24228 20700 24292 20704
rect 24228 20644 24232 20700
rect 24232 20644 24288 20700
rect 24288 20644 24292 20700
rect 24228 20640 24292 20644
rect 24308 20700 24372 20704
rect 24308 20644 24312 20700
rect 24312 20644 24368 20700
rect 24368 20644 24372 20700
rect 24308 20640 24372 20644
rect 24388 20700 24452 20704
rect 24388 20644 24392 20700
rect 24392 20644 24448 20700
rect 24448 20644 24452 20700
rect 24388 20640 24452 20644
rect 15516 20436 15580 20500
rect 4171 20156 4235 20160
rect 4171 20100 4175 20156
rect 4175 20100 4231 20156
rect 4231 20100 4235 20156
rect 4171 20096 4235 20100
rect 4251 20156 4315 20160
rect 4251 20100 4255 20156
rect 4255 20100 4311 20156
rect 4311 20100 4315 20156
rect 4251 20096 4315 20100
rect 4331 20156 4395 20160
rect 4331 20100 4335 20156
rect 4335 20100 4391 20156
rect 4391 20100 4395 20156
rect 4331 20096 4395 20100
rect 4411 20156 4475 20160
rect 4411 20100 4415 20156
rect 4415 20100 4471 20156
rect 4471 20100 4475 20156
rect 4411 20096 4475 20100
rect 10610 20156 10674 20160
rect 10610 20100 10614 20156
rect 10614 20100 10670 20156
rect 10670 20100 10674 20156
rect 10610 20096 10674 20100
rect 10690 20156 10754 20160
rect 10690 20100 10694 20156
rect 10694 20100 10750 20156
rect 10750 20100 10754 20156
rect 10690 20096 10754 20100
rect 10770 20156 10834 20160
rect 10770 20100 10774 20156
rect 10774 20100 10830 20156
rect 10830 20100 10834 20156
rect 10770 20096 10834 20100
rect 10850 20156 10914 20160
rect 10850 20100 10854 20156
rect 10854 20100 10910 20156
rect 10910 20100 10914 20156
rect 10850 20096 10914 20100
rect 17049 20156 17113 20160
rect 17049 20100 17053 20156
rect 17053 20100 17109 20156
rect 17109 20100 17113 20156
rect 17049 20096 17113 20100
rect 17129 20156 17193 20160
rect 17129 20100 17133 20156
rect 17133 20100 17189 20156
rect 17189 20100 17193 20156
rect 17129 20096 17193 20100
rect 17209 20156 17273 20160
rect 17209 20100 17213 20156
rect 17213 20100 17269 20156
rect 17269 20100 17273 20156
rect 17209 20096 17273 20100
rect 17289 20156 17353 20160
rect 17289 20100 17293 20156
rect 17293 20100 17349 20156
rect 17349 20100 17353 20156
rect 17289 20096 17353 20100
rect 23488 20156 23552 20160
rect 23488 20100 23492 20156
rect 23492 20100 23548 20156
rect 23548 20100 23552 20156
rect 23488 20096 23552 20100
rect 23568 20156 23632 20160
rect 23568 20100 23572 20156
rect 23572 20100 23628 20156
rect 23628 20100 23632 20156
rect 23568 20096 23632 20100
rect 23648 20156 23712 20160
rect 23648 20100 23652 20156
rect 23652 20100 23708 20156
rect 23708 20100 23712 20156
rect 23648 20096 23712 20100
rect 23728 20156 23792 20160
rect 23728 20100 23732 20156
rect 23732 20100 23788 20156
rect 23788 20100 23792 20156
rect 23728 20096 23792 20100
rect 4831 19612 4895 19616
rect 4831 19556 4835 19612
rect 4835 19556 4891 19612
rect 4891 19556 4895 19612
rect 4831 19552 4895 19556
rect 4911 19612 4975 19616
rect 4911 19556 4915 19612
rect 4915 19556 4971 19612
rect 4971 19556 4975 19612
rect 4911 19552 4975 19556
rect 4991 19612 5055 19616
rect 4991 19556 4995 19612
rect 4995 19556 5051 19612
rect 5051 19556 5055 19612
rect 4991 19552 5055 19556
rect 5071 19612 5135 19616
rect 5071 19556 5075 19612
rect 5075 19556 5131 19612
rect 5131 19556 5135 19612
rect 5071 19552 5135 19556
rect 11270 19612 11334 19616
rect 11270 19556 11274 19612
rect 11274 19556 11330 19612
rect 11330 19556 11334 19612
rect 11270 19552 11334 19556
rect 11350 19612 11414 19616
rect 11350 19556 11354 19612
rect 11354 19556 11410 19612
rect 11410 19556 11414 19612
rect 11350 19552 11414 19556
rect 11430 19612 11494 19616
rect 11430 19556 11434 19612
rect 11434 19556 11490 19612
rect 11490 19556 11494 19612
rect 11430 19552 11494 19556
rect 11510 19612 11574 19616
rect 11510 19556 11514 19612
rect 11514 19556 11570 19612
rect 11570 19556 11574 19612
rect 11510 19552 11574 19556
rect 17709 19612 17773 19616
rect 17709 19556 17713 19612
rect 17713 19556 17769 19612
rect 17769 19556 17773 19612
rect 17709 19552 17773 19556
rect 17789 19612 17853 19616
rect 17789 19556 17793 19612
rect 17793 19556 17849 19612
rect 17849 19556 17853 19612
rect 17789 19552 17853 19556
rect 17869 19612 17933 19616
rect 17869 19556 17873 19612
rect 17873 19556 17929 19612
rect 17929 19556 17933 19612
rect 17869 19552 17933 19556
rect 17949 19612 18013 19616
rect 17949 19556 17953 19612
rect 17953 19556 18009 19612
rect 18009 19556 18013 19612
rect 17949 19552 18013 19556
rect 24148 19612 24212 19616
rect 24148 19556 24152 19612
rect 24152 19556 24208 19612
rect 24208 19556 24212 19612
rect 24148 19552 24212 19556
rect 24228 19612 24292 19616
rect 24228 19556 24232 19612
rect 24232 19556 24288 19612
rect 24288 19556 24292 19612
rect 24228 19552 24292 19556
rect 24308 19612 24372 19616
rect 24308 19556 24312 19612
rect 24312 19556 24368 19612
rect 24368 19556 24372 19612
rect 24308 19552 24372 19556
rect 24388 19612 24452 19616
rect 24388 19556 24392 19612
rect 24392 19556 24448 19612
rect 24448 19556 24452 19612
rect 24388 19552 24452 19556
rect 4171 19068 4235 19072
rect 4171 19012 4175 19068
rect 4175 19012 4231 19068
rect 4231 19012 4235 19068
rect 4171 19008 4235 19012
rect 4251 19068 4315 19072
rect 4251 19012 4255 19068
rect 4255 19012 4311 19068
rect 4311 19012 4315 19068
rect 4251 19008 4315 19012
rect 4331 19068 4395 19072
rect 4331 19012 4335 19068
rect 4335 19012 4391 19068
rect 4391 19012 4395 19068
rect 4331 19008 4395 19012
rect 4411 19068 4475 19072
rect 4411 19012 4415 19068
rect 4415 19012 4471 19068
rect 4471 19012 4475 19068
rect 4411 19008 4475 19012
rect 10610 19068 10674 19072
rect 10610 19012 10614 19068
rect 10614 19012 10670 19068
rect 10670 19012 10674 19068
rect 10610 19008 10674 19012
rect 10690 19068 10754 19072
rect 10690 19012 10694 19068
rect 10694 19012 10750 19068
rect 10750 19012 10754 19068
rect 10690 19008 10754 19012
rect 10770 19068 10834 19072
rect 10770 19012 10774 19068
rect 10774 19012 10830 19068
rect 10830 19012 10834 19068
rect 10770 19008 10834 19012
rect 10850 19068 10914 19072
rect 10850 19012 10854 19068
rect 10854 19012 10910 19068
rect 10910 19012 10914 19068
rect 10850 19008 10914 19012
rect 17049 19068 17113 19072
rect 17049 19012 17053 19068
rect 17053 19012 17109 19068
rect 17109 19012 17113 19068
rect 17049 19008 17113 19012
rect 17129 19068 17193 19072
rect 17129 19012 17133 19068
rect 17133 19012 17189 19068
rect 17189 19012 17193 19068
rect 17129 19008 17193 19012
rect 17209 19068 17273 19072
rect 17209 19012 17213 19068
rect 17213 19012 17269 19068
rect 17269 19012 17273 19068
rect 17209 19008 17273 19012
rect 17289 19068 17353 19072
rect 17289 19012 17293 19068
rect 17293 19012 17349 19068
rect 17349 19012 17353 19068
rect 17289 19008 17353 19012
rect 23488 19068 23552 19072
rect 23488 19012 23492 19068
rect 23492 19012 23548 19068
rect 23548 19012 23552 19068
rect 23488 19008 23552 19012
rect 23568 19068 23632 19072
rect 23568 19012 23572 19068
rect 23572 19012 23628 19068
rect 23628 19012 23632 19068
rect 23568 19008 23632 19012
rect 23648 19068 23712 19072
rect 23648 19012 23652 19068
rect 23652 19012 23708 19068
rect 23708 19012 23712 19068
rect 23648 19008 23712 19012
rect 23728 19068 23792 19072
rect 23728 19012 23732 19068
rect 23732 19012 23788 19068
rect 23788 19012 23792 19068
rect 23728 19008 23792 19012
rect 4831 18524 4895 18528
rect 4831 18468 4835 18524
rect 4835 18468 4891 18524
rect 4891 18468 4895 18524
rect 4831 18464 4895 18468
rect 4911 18524 4975 18528
rect 4911 18468 4915 18524
rect 4915 18468 4971 18524
rect 4971 18468 4975 18524
rect 4911 18464 4975 18468
rect 4991 18524 5055 18528
rect 4991 18468 4995 18524
rect 4995 18468 5051 18524
rect 5051 18468 5055 18524
rect 4991 18464 5055 18468
rect 5071 18524 5135 18528
rect 5071 18468 5075 18524
rect 5075 18468 5131 18524
rect 5131 18468 5135 18524
rect 5071 18464 5135 18468
rect 11270 18524 11334 18528
rect 11270 18468 11274 18524
rect 11274 18468 11330 18524
rect 11330 18468 11334 18524
rect 11270 18464 11334 18468
rect 11350 18524 11414 18528
rect 11350 18468 11354 18524
rect 11354 18468 11410 18524
rect 11410 18468 11414 18524
rect 11350 18464 11414 18468
rect 11430 18524 11494 18528
rect 11430 18468 11434 18524
rect 11434 18468 11490 18524
rect 11490 18468 11494 18524
rect 11430 18464 11494 18468
rect 11510 18524 11574 18528
rect 11510 18468 11514 18524
rect 11514 18468 11570 18524
rect 11570 18468 11574 18524
rect 11510 18464 11574 18468
rect 17709 18524 17773 18528
rect 17709 18468 17713 18524
rect 17713 18468 17769 18524
rect 17769 18468 17773 18524
rect 17709 18464 17773 18468
rect 17789 18524 17853 18528
rect 17789 18468 17793 18524
rect 17793 18468 17849 18524
rect 17849 18468 17853 18524
rect 17789 18464 17853 18468
rect 17869 18524 17933 18528
rect 17869 18468 17873 18524
rect 17873 18468 17929 18524
rect 17929 18468 17933 18524
rect 17869 18464 17933 18468
rect 17949 18524 18013 18528
rect 17949 18468 17953 18524
rect 17953 18468 18009 18524
rect 18009 18468 18013 18524
rect 17949 18464 18013 18468
rect 24148 18524 24212 18528
rect 24148 18468 24152 18524
rect 24152 18468 24208 18524
rect 24208 18468 24212 18524
rect 24148 18464 24212 18468
rect 24228 18524 24292 18528
rect 24228 18468 24232 18524
rect 24232 18468 24288 18524
rect 24288 18468 24292 18524
rect 24228 18464 24292 18468
rect 24308 18524 24372 18528
rect 24308 18468 24312 18524
rect 24312 18468 24368 18524
rect 24368 18468 24372 18524
rect 24308 18464 24372 18468
rect 24388 18524 24452 18528
rect 24388 18468 24392 18524
rect 24392 18468 24448 18524
rect 24448 18468 24452 18524
rect 24388 18464 24452 18468
rect 4171 17980 4235 17984
rect 4171 17924 4175 17980
rect 4175 17924 4231 17980
rect 4231 17924 4235 17980
rect 4171 17920 4235 17924
rect 4251 17980 4315 17984
rect 4251 17924 4255 17980
rect 4255 17924 4311 17980
rect 4311 17924 4315 17980
rect 4251 17920 4315 17924
rect 4331 17980 4395 17984
rect 4331 17924 4335 17980
rect 4335 17924 4391 17980
rect 4391 17924 4395 17980
rect 4331 17920 4395 17924
rect 4411 17980 4475 17984
rect 4411 17924 4415 17980
rect 4415 17924 4471 17980
rect 4471 17924 4475 17980
rect 4411 17920 4475 17924
rect 10610 17980 10674 17984
rect 10610 17924 10614 17980
rect 10614 17924 10670 17980
rect 10670 17924 10674 17980
rect 10610 17920 10674 17924
rect 10690 17980 10754 17984
rect 10690 17924 10694 17980
rect 10694 17924 10750 17980
rect 10750 17924 10754 17980
rect 10690 17920 10754 17924
rect 10770 17980 10834 17984
rect 10770 17924 10774 17980
rect 10774 17924 10830 17980
rect 10830 17924 10834 17980
rect 10770 17920 10834 17924
rect 10850 17980 10914 17984
rect 10850 17924 10854 17980
rect 10854 17924 10910 17980
rect 10910 17924 10914 17980
rect 10850 17920 10914 17924
rect 17049 17980 17113 17984
rect 17049 17924 17053 17980
rect 17053 17924 17109 17980
rect 17109 17924 17113 17980
rect 17049 17920 17113 17924
rect 17129 17980 17193 17984
rect 17129 17924 17133 17980
rect 17133 17924 17189 17980
rect 17189 17924 17193 17980
rect 17129 17920 17193 17924
rect 17209 17980 17273 17984
rect 17209 17924 17213 17980
rect 17213 17924 17269 17980
rect 17269 17924 17273 17980
rect 17209 17920 17273 17924
rect 17289 17980 17353 17984
rect 17289 17924 17293 17980
rect 17293 17924 17349 17980
rect 17349 17924 17353 17980
rect 17289 17920 17353 17924
rect 23488 17980 23552 17984
rect 23488 17924 23492 17980
rect 23492 17924 23548 17980
rect 23548 17924 23552 17980
rect 23488 17920 23552 17924
rect 23568 17980 23632 17984
rect 23568 17924 23572 17980
rect 23572 17924 23628 17980
rect 23628 17924 23632 17980
rect 23568 17920 23632 17924
rect 23648 17980 23712 17984
rect 23648 17924 23652 17980
rect 23652 17924 23708 17980
rect 23708 17924 23712 17980
rect 23648 17920 23712 17924
rect 23728 17980 23792 17984
rect 23728 17924 23732 17980
rect 23732 17924 23788 17980
rect 23788 17924 23792 17980
rect 23728 17920 23792 17924
rect 15516 17912 15580 17916
rect 15516 17856 15530 17912
rect 15530 17856 15580 17912
rect 15516 17852 15580 17856
rect 4831 17436 4895 17440
rect 4831 17380 4835 17436
rect 4835 17380 4891 17436
rect 4891 17380 4895 17436
rect 4831 17376 4895 17380
rect 4911 17436 4975 17440
rect 4911 17380 4915 17436
rect 4915 17380 4971 17436
rect 4971 17380 4975 17436
rect 4911 17376 4975 17380
rect 4991 17436 5055 17440
rect 4991 17380 4995 17436
rect 4995 17380 5051 17436
rect 5051 17380 5055 17436
rect 4991 17376 5055 17380
rect 5071 17436 5135 17440
rect 5071 17380 5075 17436
rect 5075 17380 5131 17436
rect 5131 17380 5135 17436
rect 5071 17376 5135 17380
rect 11270 17436 11334 17440
rect 11270 17380 11274 17436
rect 11274 17380 11330 17436
rect 11330 17380 11334 17436
rect 11270 17376 11334 17380
rect 11350 17436 11414 17440
rect 11350 17380 11354 17436
rect 11354 17380 11410 17436
rect 11410 17380 11414 17436
rect 11350 17376 11414 17380
rect 11430 17436 11494 17440
rect 11430 17380 11434 17436
rect 11434 17380 11490 17436
rect 11490 17380 11494 17436
rect 11430 17376 11494 17380
rect 11510 17436 11574 17440
rect 11510 17380 11514 17436
rect 11514 17380 11570 17436
rect 11570 17380 11574 17436
rect 11510 17376 11574 17380
rect 17709 17436 17773 17440
rect 17709 17380 17713 17436
rect 17713 17380 17769 17436
rect 17769 17380 17773 17436
rect 17709 17376 17773 17380
rect 17789 17436 17853 17440
rect 17789 17380 17793 17436
rect 17793 17380 17849 17436
rect 17849 17380 17853 17436
rect 17789 17376 17853 17380
rect 17869 17436 17933 17440
rect 17869 17380 17873 17436
rect 17873 17380 17929 17436
rect 17929 17380 17933 17436
rect 17869 17376 17933 17380
rect 17949 17436 18013 17440
rect 17949 17380 17953 17436
rect 17953 17380 18009 17436
rect 18009 17380 18013 17436
rect 17949 17376 18013 17380
rect 24148 17436 24212 17440
rect 24148 17380 24152 17436
rect 24152 17380 24208 17436
rect 24208 17380 24212 17436
rect 24148 17376 24212 17380
rect 24228 17436 24292 17440
rect 24228 17380 24232 17436
rect 24232 17380 24288 17436
rect 24288 17380 24292 17436
rect 24228 17376 24292 17380
rect 24308 17436 24372 17440
rect 24308 17380 24312 17436
rect 24312 17380 24368 17436
rect 24368 17380 24372 17436
rect 24308 17376 24372 17380
rect 24388 17436 24452 17440
rect 24388 17380 24392 17436
rect 24392 17380 24448 17436
rect 24448 17380 24452 17436
rect 24388 17376 24452 17380
rect 15332 17368 15396 17372
rect 15332 17312 15382 17368
rect 15382 17312 15396 17368
rect 15332 17308 15396 17312
rect 4171 16892 4235 16896
rect 4171 16836 4175 16892
rect 4175 16836 4231 16892
rect 4231 16836 4235 16892
rect 4171 16832 4235 16836
rect 4251 16892 4315 16896
rect 4251 16836 4255 16892
rect 4255 16836 4311 16892
rect 4311 16836 4315 16892
rect 4251 16832 4315 16836
rect 4331 16892 4395 16896
rect 4331 16836 4335 16892
rect 4335 16836 4391 16892
rect 4391 16836 4395 16892
rect 4331 16832 4395 16836
rect 4411 16892 4475 16896
rect 4411 16836 4415 16892
rect 4415 16836 4471 16892
rect 4471 16836 4475 16892
rect 4411 16832 4475 16836
rect 10610 16892 10674 16896
rect 10610 16836 10614 16892
rect 10614 16836 10670 16892
rect 10670 16836 10674 16892
rect 10610 16832 10674 16836
rect 10690 16892 10754 16896
rect 10690 16836 10694 16892
rect 10694 16836 10750 16892
rect 10750 16836 10754 16892
rect 10690 16832 10754 16836
rect 10770 16892 10834 16896
rect 10770 16836 10774 16892
rect 10774 16836 10830 16892
rect 10830 16836 10834 16892
rect 10770 16832 10834 16836
rect 10850 16892 10914 16896
rect 10850 16836 10854 16892
rect 10854 16836 10910 16892
rect 10910 16836 10914 16892
rect 10850 16832 10914 16836
rect 17049 16892 17113 16896
rect 17049 16836 17053 16892
rect 17053 16836 17109 16892
rect 17109 16836 17113 16892
rect 17049 16832 17113 16836
rect 17129 16892 17193 16896
rect 17129 16836 17133 16892
rect 17133 16836 17189 16892
rect 17189 16836 17193 16892
rect 17129 16832 17193 16836
rect 17209 16892 17273 16896
rect 17209 16836 17213 16892
rect 17213 16836 17269 16892
rect 17269 16836 17273 16892
rect 17209 16832 17273 16836
rect 17289 16892 17353 16896
rect 17289 16836 17293 16892
rect 17293 16836 17349 16892
rect 17349 16836 17353 16892
rect 17289 16832 17353 16836
rect 23488 16892 23552 16896
rect 23488 16836 23492 16892
rect 23492 16836 23548 16892
rect 23548 16836 23552 16892
rect 23488 16832 23552 16836
rect 23568 16892 23632 16896
rect 23568 16836 23572 16892
rect 23572 16836 23628 16892
rect 23628 16836 23632 16892
rect 23568 16832 23632 16836
rect 23648 16892 23712 16896
rect 23648 16836 23652 16892
rect 23652 16836 23708 16892
rect 23708 16836 23712 16892
rect 23648 16832 23712 16836
rect 23728 16892 23792 16896
rect 23728 16836 23732 16892
rect 23732 16836 23788 16892
rect 23788 16836 23792 16892
rect 23728 16832 23792 16836
rect 4831 16348 4895 16352
rect 4831 16292 4835 16348
rect 4835 16292 4891 16348
rect 4891 16292 4895 16348
rect 4831 16288 4895 16292
rect 4911 16348 4975 16352
rect 4911 16292 4915 16348
rect 4915 16292 4971 16348
rect 4971 16292 4975 16348
rect 4911 16288 4975 16292
rect 4991 16348 5055 16352
rect 4991 16292 4995 16348
rect 4995 16292 5051 16348
rect 5051 16292 5055 16348
rect 4991 16288 5055 16292
rect 5071 16348 5135 16352
rect 5071 16292 5075 16348
rect 5075 16292 5131 16348
rect 5131 16292 5135 16348
rect 5071 16288 5135 16292
rect 11270 16348 11334 16352
rect 11270 16292 11274 16348
rect 11274 16292 11330 16348
rect 11330 16292 11334 16348
rect 11270 16288 11334 16292
rect 11350 16348 11414 16352
rect 11350 16292 11354 16348
rect 11354 16292 11410 16348
rect 11410 16292 11414 16348
rect 11350 16288 11414 16292
rect 11430 16348 11494 16352
rect 11430 16292 11434 16348
rect 11434 16292 11490 16348
rect 11490 16292 11494 16348
rect 11430 16288 11494 16292
rect 11510 16348 11574 16352
rect 11510 16292 11514 16348
rect 11514 16292 11570 16348
rect 11570 16292 11574 16348
rect 11510 16288 11574 16292
rect 17709 16348 17773 16352
rect 17709 16292 17713 16348
rect 17713 16292 17769 16348
rect 17769 16292 17773 16348
rect 17709 16288 17773 16292
rect 17789 16348 17853 16352
rect 17789 16292 17793 16348
rect 17793 16292 17849 16348
rect 17849 16292 17853 16348
rect 17789 16288 17853 16292
rect 17869 16348 17933 16352
rect 17869 16292 17873 16348
rect 17873 16292 17929 16348
rect 17929 16292 17933 16348
rect 17869 16288 17933 16292
rect 17949 16348 18013 16352
rect 17949 16292 17953 16348
rect 17953 16292 18009 16348
rect 18009 16292 18013 16348
rect 17949 16288 18013 16292
rect 24148 16348 24212 16352
rect 24148 16292 24152 16348
rect 24152 16292 24208 16348
rect 24208 16292 24212 16348
rect 24148 16288 24212 16292
rect 24228 16348 24292 16352
rect 24228 16292 24232 16348
rect 24232 16292 24288 16348
rect 24288 16292 24292 16348
rect 24228 16288 24292 16292
rect 24308 16348 24372 16352
rect 24308 16292 24312 16348
rect 24312 16292 24368 16348
rect 24368 16292 24372 16348
rect 24308 16288 24372 16292
rect 24388 16348 24452 16352
rect 24388 16292 24392 16348
rect 24392 16292 24448 16348
rect 24448 16292 24452 16348
rect 24388 16288 24452 16292
rect 4171 15804 4235 15808
rect 4171 15748 4175 15804
rect 4175 15748 4231 15804
rect 4231 15748 4235 15804
rect 4171 15744 4235 15748
rect 4251 15804 4315 15808
rect 4251 15748 4255 15804
rect 4255 15748 4311 15804
rect 4311 15748 4315 15804
rect 4251 15744 4315 15748
rect 4331 15804 4395 15808
rect 4331 15748 4335 15804
rect 4335 15748 4391 15804
rect 4391 15748 4395 15804
rect 4331 15744 4395 15748
rect 4411 15804 4475 15808
rect 4411 15748 4415 15804
rect 4415 15748 4471 15804
rect 4471 15748 4475 15804
rect 4411 15744 4475 15748
rect 10610 15804 10674 15808
rect 10610 15748 10614 15804
rect 10614 15748 10670 15804
rect 10670 15748 10674 15804
rect 10610 15744 10674 15748
rect 10690 15804 10754 15808
rect 10690 15748 10694 15804
rect 10694 15748 10750 15804
rect 10750 15748 10754 15804
rect 10690 15744 10754 15748
rect 10770 15804 10834 15808
rect 10770 15748 10774 15804
rect 10774 15748 10830 15804
rect 10830 15748 10834 15804
rect 10770 15744 10834 15748
rect 10850 15804 10914 15808
rect 10850 15748 10854 15804
rect 10854 15748 10910 15804
rect 10910 15748 10914 15804
rect 10850 15744 10914 15748
rect 17049 15804 17113 15808
rect 17049 15748 17053 15804
rect 17053 15748 17109 15804
rect 17109 15748 17113 15804
rect 17049 15744 17113 15748
rect 17129 15804 17193 15808
rect 17129 15748 17133 15804
rect 17133 15748 17189 15804
rect 17189 15748 17193 15804
rect 17129 15744 17193 15748
rect 17209 15804 17273 15808
rect 17209 15748 17213 15804
rect 17213 15748 17269 15804
rect 17269 15748 17273 15804
rect 17209 15744 17273 15748
rect 17289 15804 17353 15808
rect 17289 15748 17293 15804
rect 17293 15748 17349 15804
rect 17349 15748 17353 15804
rect 17289 15744 17353 15748
rect 23488 15804 23552 15808
rect 23488 15748 23492 15804
rect 23492 15748 23548 15804
rect 23548 15748 23552 15804
rect 23488 15744 23552 15748
rect 23568 15804 23632 15808
rect 23568 15748 23572 15804
rect 23572 15748 23628 15804
rect 23628 15748 23632 15804
rect 23568 15744 23632 15748
rect 23648 15804 23712 15808
rect 23648 15748 23652 15804
rect 23652 15748 23708 15804
rect 23708 15748 23712 15804
rect 23648 15744 23712 15748
rect 23728 15804 23792 15808
rect 23728 15748 23732 15804
rect 23732 15748 23788 15804
rect 23788 15748 23792 15804
rect 23728 15744 23792 15748
rect 4831 15260 4895 15264
rect 4831 15204 4835 15260
rect 4835 15204 4891 15260
rect 4891 15204 4895 15260
rect 4831 15200 4895 15204
rect 4911 15260 4975 15264
rect 4911 15204 4915 15260
rect 4915 15204 4971 15260
rect 4971 15204 4975 15260
rect 4911 15200 4975 15204
rect 4991 15260 5055 15264
rect 4991 15204 4995 15260
rect 4995 15204 5051 15260
rect 5051 15204 5055 15260
rect 4991 15200 5055 15204
rect 5071 15260 5135 15264
rect 5071 15204 5075 15260
rect 5075 15204 5131 15260
rect 5131 15204 5135 15260
rect 5071 15200 5135 15204
rect 11270 15260 11334 15264
rect 11270 15204 11274 15260
rect 11274 15204 11330 15260
rect 11330 15204 11334 15260
rect 11270 15200 11334 15204
rect 11350 15260 11414 15264
rect 11350 15204 11354 15260
rect 11354 15204 11410 15260
rect 11410 15204 11414 15260
rect 11350 15200 11414 15204
rect 11430 15260 11494 15264
rect 11430 15204 11434 15260
rect 11434 15204 11490 15260
rect 11490 15204 11494 15260
rect 11430 15200 11494 15204
rect 11510 15260 11574 15264
rect 11510 15204 11514 15260
rect 11514 15204 11570 15260
rect 11570 15204 11574 15260
rect 11510 15200 11574 15204
rect 17709 15260 17773 15264
rect 17709 15204 17713 15260
rect 17713 15204 17769 15260
rect 17769 15204 17773 15260
rect 17709 15200 17773 15204
rect 17789 15260 17853 15264
rect 17789 15204 17793 15260
rect 17793 15204 17849 15260
rect 17849 15204 17853 15260
rect 17789 15200 17853 15204
rect 17869 15260 17933 15264
rect 17869 15204 17873 15260
rect 17873 15204 17929 15260
rect 17929 15204 17933 15260
rect 17869 15200 17933 15204
rect 17949 15260 18013 15264
rect 17949 15204 17953 15260
rect 17953 15204 18009 15260
rect 18009 15204 18013 15260
rect 17949 15200 18013 15204
rect 24148 15260 24212 15264
rect 24148 15204 24152 15260
rect 24152 15204 24208 15260
rect 24208 15204 24212 15260
rect 24148 15200 24212 15204
rect 24228 15260 24292 15264
rect 24228 15204 24232 15260
rect 24232 15204 24288 15260
rect 24288 15204 24292 15260
rect 24228 15200 24292 15204
rect 24308 15260 24372 15264
rect 24308 15204 24312 15260
rect 24312 15204 24368 15260
rect 24368 15204 24372 15260
rect 24308 15200 24372 15204
rect 24388 15260 24452 15264
rect 24388 15204 24392 15260
rect 24392 15204 24448 15260
rect 24448 15204 24452 15260
rect 24388 15200 24452 15204
rect 4171 14716 4235 14720
rect 4171 14660 4175 14716
rect 4175 14660 4231 14716
rect 4231 14660 4235 14716
rect 4171 14656 4235 14660
rect 4251 14716 4315 14720
rect 4251 14660 4255 14716
rect 4255 14660 4311 14716
rect 4311 14660 4315 14716
rect 4251 14656 4315 14660
rect 4331 14716 4395 14720
rect 4331 14660 4335 14716
rect 4335 14660 4391 14716
rect 4391 14660 4395 14716
rect 4331 14656 4395 14660
rect 4411 14716 4475 14720
rect 4411 14660 4415 14716
rect 4415 14660 4471 14716
rect 4471 14660 4475 14716
rect 4411 14656 4475 14660
rect 10610 14716 10674 14720
rect 10610 14660 10614 14716
rect 10614 14660 10670 14716
rect 10670 14660 10674 14716
rect 10610 14656 10674 14660
rect 10690 14716 10754 14720
rect 10690 14660 10694 14716
rect 10694 14660 10750 14716
rect 10750 14660 10754 14716
rect 10690 14656 10754 14660
rect 10770 14716 10834 14720
rect 10770 14660 10774 14716
rect 10774 14660 10830 14716
rect 10830 14660 10834 14716
rect 10770 14656 10834 14660
rect 10850 14716 10914 14720
rect 10850 14660 10854 14716
rect 10854 14660 10910 14716
rect 10910 14660 10914 14716
rect 10850 14656 10914 14660
rect 17049 14716 17113 14720
rect 17049 14660 17053 14716
rect 17053 14660 17109 14716
rect 17109 14660 17113 14716
rect 17049 14656 17113 14660
rect 17129 14716 17193 14720
rect 17129 14660 17133 14716
rect 17133 14660 17189 14716
rect 17189 14660 17193 14716
rect 17129 14656 17193 14660
rect 17209 14716 17273 14720
rect 17209 14660 17213 14716
rect 17213 14660 17269 14716
rect 17269 14660 17273 14716
rect 17209 14656 17273 14660
rect 17289 14716 17353 14720
rect 17289 14660 17293 14716
rect 17293 14660 17349 14716
rect 17349 14660 17353 14716
rect 17289 14656 17353 14660
rect 23488 14716 23552 14720
rect 23488 14660 23492 14716
rect 23492 14660 23548 14716
rect 23548 14660 23552 14716
rect 23488 14656 23552 14660
rect 23568 14716 23632 14720
rect 23568 14660 23572 14716
rect 23572 14660 23628 14716
rect 23628 14660 23632 14716
rect 23568 14656 23632 14660
rect 23648 14716 23712 14720
rect 23648 14660 23652 14716
rect 23652 14660 23708 14716
rect 23708 14660 23712 14716
rect 23648 14656 23712 14660
rect 23728 14716 23792 14720
rect 23728 14660 23732 14716
rect 23732 14660 23788 14716
rect 23788 14660 23792 14716
rect 23728 14656 23792 14660
rect 4831 14172 4895 14176
rect 4831 14116 4835 14172
rect 4835 14116 4891 14172
rect 4891 14116 4895 14172
rect 4831 14112 4895 14116
rect 4911 14172 4975 14176
rect 4911 14116 4915 14172
rect 4915 14116 4971 14172
rect 4971 14116 4975 14172
rect 4911 14112 4975 14116
rect 4991 14172 5055 14176
rect 4991 14116 4995 14172
rect 4995 14116 5051 14172
rect 5051 14116 5055 14172
rect 4991 14112 5055 14116
rect 5071 14172 5135 14176
rect 5071 14116 5075 14172
rect 5075 14116 5131 14172
rect 5131 14116 5135 14172
rect 5071 14112 5135 14116
rect 11270 14172 11334 14176
rect 11270 14116 11274 14172
rect 11274 14116 11330 14172
rect 11330 14116 11334 14172
rect 11270 14112 11334 14116
rect 11350 14172 11414 14176
rect 11350 14116 11354 14172
rect 11354 14116 11410 14172
rect 11410 14116 11414 14172
rect 11350 14112 11414 14116
rect 11430 14172 11494 14176
rect 11430 14116 11434 14172
rect 11434 14116 11490 14172
rect 11490 14116 11494 14172
rect 11430 14112 11494 14116
rect 11510 14172 11574 14176
rect 11510 14116 11514 14172
rect 11514 14116 11570 14172
rect 11570 14116 11574 14172
rect 11510 14112 11574 14116
rect 17709 14172 17773 14176
rect 17709 14116 17713 14172
rect 17713 14116 17769 14172
rect 17769 14116 17773 14172
rect 17709 14112 17773 14116
rect 17789 14172 17853 14176
rect 17789 14116 17793 14172
rect 17793 14116 17849 14172
rect 17849 14116 17853 14172
rect 17789 14112 17853 14116
rect 17869 14172 17933 14176
rect 17869 14116 17873 14172
rect 17873 14116 17929 14172
rect 17929 14116 17933 14172
rect 17869 14112 17933 14116
rect 17949 14172 18013 14176
rect 17949 14116 17953 14172
rect 17953 14116 18009 14172
rect 18009 14116 18013 14172
rect 17949 14112 18013 14116
rect 24148 14172 24212 14176
rect 24148 14116 24152 14172
rect 24152 14116 24208 14172
rect 24208 14116 24212 14172
rect 24148 14112 24212 14116
rect 24228 14172 24292 14176
rect 24228 14116 24232 14172
rect 24232 14116 24288 14172
rect 24288 14116 24292 14172
rect 24228 14112 24292 14116
rect 24308 14172 24372 14176
rect 24308 14116 24312 14172
rect 24312 14116 24368 14172
rect 24368 14116 24372 14172
rect 24308 14112 24372 14116
rect 24388 14172 24452 14176
rect 24388 14116 24392 14172
rect 24392 14116 24448 14172
rect 24448 14116 24452 14172
rect 24388 14112 24452 14116
rect 4171 13628 4235 13632
rect 4171 13572 4175 13628
rect 4175 13572 4231 13628
rect 4231 13572 4235 13628
rect 4171 13568 4235 13572
rect 4251 13628 4315 13632
rect 4251 13572 4255 13628
rect 4255 13572 4311 13628
rect 4311 13572 4315 13628
rect 4251 13568 4315 13572
rect 4331 13628 4395 13632
rect 4331 13572 4335 13628
rect 4335 13572 4391 13628
rect 4391 13572 4395 13628
rect 4331 13568 4395 13572
rect 4411 13628 4475 13632
rect 4411 13572 4415 13628
rect 4415 13572 4471 13628
rect 4471 13572 4475 13628
rect 4411 13568 4475 13572
rect 10610 13628 10674 13632
rect 10610 13572 10614 13628
rect 10614 13572 10670 13628
rect 10670 13572 10674 13628
rect 10610 13568 10674 13572
rect 10690 13628 10754 13632
rect 10690 13572 10694 13628
rect 10694 13572 10750 13628
rect 10750 13572 10754 13628
rect 10690 13568 10754 13572
rect 10770 13628 10834 13632
rect 10770 13572 10774 13628
rect 10774 13572 10830 13628
rect 10830 13572 10834 13628
rect 10770 13568 10834 13572
rect 10850 13628 10914 13632
rect 10850 13572 10854 13628
rect 10854 13572 10910 13628
rect 10910 13572 10914 13628
rect 10850 13568 10914 13572
rect 17049 13628 17113 13632
rect 17049 13572 17053 13628
rect 17053 13572 17109 13628
rect 17109 13572 17113 13628
rect 17049 13568 17113 13572
rect 17129 13628 17193 13632
rect 17129 13572 17133 13628
rect 17133 13572 17189 13628
rect 17189 13572 17193 13628
rect 17129 13568 17193 13572
rect 17209 13628 17273 13632
rect 17209 13572 17213 13628
rect 17213 13572 17269 13628
rect 17269 13572 17273 13628
rect 17209 13568 17273 13572
rect 17289 13628 17353 13632
rect 17289 13572 17293 13628
rect 17293 13572 17349 13628
rect 17349 13572 17353 13628
rect 17289 13568 17353 13572
rect 23488 13628 23552 13632
rect 23488 13572 23492 13628
rect 23492 13572 23548 13628
rect 23548 13572 23552 13628
rect 23488 13568 23552 13572
rect 23568 13628 23632 13632
rect 23568 13572 23572 13628
rect 23572 13572 23628 13628
rect 23628 13572 23632 13628
rect 23568 13568 23632 13572
rect 23648 13628 23712 13632
rect 23648 13572 23652 13628
rect 23652 13572 23708 13628
rect 23708 13572 23712 13628
rect 23648 13568 23712 13572
rect 23728 13628 23792 13632
rect 23728 13572 23732 13628
rect 23732 13572 23788 13628
rect 23788 13572 23792 13628
rect 23728 13568 23792 13572
rect 4831 13084 4895 13088
rect 4831 13028 4835 13084
rect 4835 13028 4891 13084
rect 4891 13028 4895 13084
rect 4831 13024 4895 13028
rect 4911 13084 4975 13088
rect 4911 13028 4915 13084
rect 4915 13028 4971 13084
rect 4971 13028 4975 13084
rect 4911 13024 4975 13028
rect 4991 13084 5055 13088
rect 4991 13028 4995 13084
rect 4995 13028 5051 13084
rect 5051 13028 5055 13084
rect 4991 13024 5055 13028
rect 5071 13084 5135 13088
rect 5071 13028 5075 13084
rect 5075 13028 5131 13084
rect 5131 13028 5135 13084
rect 5071 13024 5135 13028
rect 11270 13084 11334 13088
rect 11270 13028 11274 13084
rect 11274 13028 11330 13084
rect 11330 13028 11334 13084
rect 11270 13024 11334 13028
rect 11350 13084 11414 13088
rect 11350 13028 11354 13084
rect 11354 13028 11410 13084
rect 11410 13028 11414 13084
rect 11350 13024 11414 13028
rect 11430 13084 11494 13088
rect 11430 13028 11434 13084
rect 11434 13028 11490 13084
rect 11490 13028 11494 13084
rect 11430 13024 11494 13028
rect 11510 13084 11574 13088
rect 11510 13028 11514 13084
rect 11514 13028 11570 13084
rect 11570 13028 11574 13084
rect 11510 13024 11574 13028
rect 17709 13084 17773 13088
rect 17709 13028 17713 13084
rect 17713 13028 17769 13084
rect 17769 13028 17773 13084
rect 17709 13024 17773 13028
rect 17789 13084 17853 13088
rect 17789 13028 17793 13084
rect 17793 13028 17849 13084
rect 17849 13028 17853 13084
rect 17789 13024 17853 13028
rect 17869 13084 17933 13088
rect 17869 13028 17873 13084
rect 17873 13028 17929 13084
rect 17929 13028 17933 13084
rect 17869 13024 17933 13028
rect 17949 13084 18013 13088
rect 17949 13028 17953 13084
rect 17953 13028 18009 13084
rect 18009 13028 18013 13084
rect 17949 13024 18013 13028
rect 24148 13084 24212 13088
rect 24148 13028 24152 13084
rect 24152 13028 24208 13084
rect 24208 13028 24212 13084
rect 24148 13024 24212 13028
rect 24228 13084 24292 13088
rect 24228 13028 24232 13084
rect 24232 13028 24288 13084
rect 24288 13028 24292 13084
rect 24228 13024 24292 13028
rect 24308 13084 24372 13088
rect 24308 13028 24312 13084
rect 24312 13028 24368 13084
rect 24368 13028 24372 13084
rect 24308 13024 24372 13028
rect 24388 13084 24452 13088
rect 24388 13028 24392 13084
rect 24392 13028 24448 13084
rect 24448 13028 24452 13084
rect 24388 13024 24452 13028
rect 4171 12540 4235 12544
rect 4171 12484 4175 12540
rect 4175 12484 4231 12540
rect 4231 12484 4235 12540
rect 4171 12480 4235 12484
rect 4251 12540 4315 12544
rect 4251 12484 4255 12540
rect 4255 12484 4311 12540
rect 4311 12484 4315 12540
rect 4251 12480 4315 12484
rect 4331 12540 4395 12544
rect 4331 12484 4335 12540
rect 4335 12484 4391 12540
rect 4391 12484 4395 12540
rect 4331 12480 4395 12484
rect 4411 12540 4475 12544
rect 4411 12484 4415 12540
rect 4415 12484 4471 12540
rect 4471 12484 4475 12540
rect 4411 12480 4475 12484
rect 10610 12540 10674 12544
rect 10610 12484 10614 12540
rect 10614 12484 10670 12540
rect 10670 12484 10674 12540
rect 10610 12480 10674 12484
rect 10690 12540 10754 12544
rect 10690 12484 10694 12540
rect 10694 12484 10750 12540
rect 10750 12484 10754 12540
rect 10690 12480 10754 12484
rect 10770 12540 10834 12544
rect 10770 12484 10774 12540
rect 10774 12484 10830 12540
rect 10830 12484 10834 12540
rect 10770 12480 10834 12484
rect 10850 12540 10914 12544
rect 10850 12484 10854 12540
rect 10854 12484 10910 12540
rect 10910 12484 10914 12540
rect 10850 12480 10914 12484
rect 17049 12540 17113 12544
rect 17049 12484 17053 12540
rect 17053 12484 17109 12540
rect 17109 12484 17113 12540
rect 17049 12480 17113 12484
rect 17129 12540 17193 12544
rect 17129 12484 17133 12540
rect 17133 12484 17189 12540
rect 17189 12484 17193 12540
rect 17129 12480 17193 12484
rect 17209 12540 17273 12544
rect 17209 12484 17213 12540
rect 17213 12484 17269 12540
rect 17269 12484 17273 12540
rect 17209 12480 17273 12484
rect 17289 12540 17353 12544
rect 17289 12484 17293 12540
rect 17293 12484 17349 12540
rect 17349 12484 17353 12540
rect 17289 12480 17353 12484
rect 23488 12540 23552 12544
rect 23488 12484 23492 12540
rect 23492 12484 23548 12540
rect 23548 12484 23552 12540
rect 23488 12480 23552 12484
rect 23568 12540 23632 12544
rect 23568 12484 23572 12540
rect 23572 12484 23628 12540
rect 23628 12484 23632 12540
rect 23568 12480 23632 12484
rect 23648 12540 23712 12544
rect 23648 12484 23652 12540
rect 23652 12484 23708 12540
rect 23708 12484 23712 12540
rect 23648 12480 23712 12484
rect 23728 12540 23792 12544
rect 23728 12484 23732 12540
rect 23732 12484 23788 12540
rect 23788 12484 23792 12540
rect 23728 12480 23792 12484
rect 4831 11996 4895 12000
rect 4831 11940 4835 11996
rect 4835 11940 4891 11996
rect 4891 11940 4895 11996
rect 4831 11936 4895 11940
rect 4911 11996 4975 12000
rect 4911 11940 4915 11996
rect 4915 11940 4971 11996
rect 4971 11940 4975 11996
rect 4911 11936 4975 11940
rect 4991 11996 5055 12000
rect 4991 11940 4995 11996
rect 4995 11940 5051 11996
rect 5051 11940 5055 11996
rect 4991 11936 5055 11940
rect 5071 11996 5135 12000
rect 5071 11940 5075 11996
rect 5075 11940 5131 11996
rect 5131 11940 5135 11996
rect 5071 11936 5135 11940
rect 11270 11996 11334 12000
rect 11270 11940 11274 11996
rect 11274 11940 11330 11996
rect 11330 11940 11334 11996
rect 11270 11936 11334 11940
rect 11350 11996 11414 12000
rect 11350 11940 11354 11996
rect 11354 11940 11410 11996
rect 11410 11940 11414 11996
rect 11350 11936 11414 11940
rect 11430 11996 11494 12000
rect 11430 11940 11434 11996
rect 11434 11940 11490 11996
rect 11490 11940 11494 11996
rect 11430 11936 11494 11940
rect 11510 11996 11574 12000
rect 11510 11940 11514 11996
rect 11514 11940 11570 11996
rect 11570 11940 11574 11996
rect 11510 11936 11574 11940
rect 17709 11996 17773 12000
rect 17709 11940 17713 11996
rect 17713 11940 17769 11996
rect 17769 11940 17773 11996
rect 17709 11936 17773 11940
rect 17789 11996 17853 12000
rect 17789 11940 17793 11996
rect 17793 11940 17849 11996
rect 17849 11940 17853 11996
rect 17789 11936 17853 11940
rect 17869 11996 17933 12000
rect 17869 11940 17873 11996
rect 17873 11940 17929 11996
rect 17929 11940 17933 11996
rect 17869 11936 17933 11940
rect 17949 11996 18013 12000
rect 17949 11940 17953 11996
rect 17953 11940 18009 11996
rect 18009 11940 18013 11996
rect 17949 11936 18013 11940
rect 24148 11996 24212 12000
rect 24148 11940 24152 11996
rect 24152 11940 24208 11996
rect 24208 11940 24212 11996
rect 24148 11936 24212 11940
rect 24228 11996 24292 12000
rect 24228 11940 24232 11996
rect 24232 11940 24288 11996
rect 24288 11940 24292 11996
rect 24228 11936 24292 11940
rect 24308 11996 24372 12000
rect 24308 11940 24312 11996
rect 24312 11940 24368 11996
rect 24368 11940 24372 11996
rect 24308 11936 24372 11940
rect 24388 11996 24452 12000
rect 24388 11940 24392 11996
rect 24392 11940 24448 11996
rect 24448 11940 24452 11996
rect 24388 11936 24452 11940
rect 4171 11452 4235 11456
rect 4171 11396 4175 11452
rect 4175 11396 4231 11452
rect 4231 11396 4235 11452
rect 4171 11392 4235 11396
rect 4251 11452 4315 11456
rect 4251 11396 4255 11452
rect 4255 11396 4311 11452
rect 4311 11396 4315 11452
rect 4251 11392 4315 11396
rect 4331 11452 4395 11456
rect 4331 11396 4335 11452
rect 4335 11396 4391 11452
rect 4391 11396 4395 11452
rect 4331 11392 4395 11396
rect 4411 11452 4475 11456
rect 4411 11396 4415 11452
rect 4415 11396 4471 11452
rect 4471 11396 4475 11452
rect 4411 11392 4475 11396
rect 10610 11452 10674 11456
rect 10610 11396 10614 11452
rect 10614 11396 10670 11452
rect 10670 11396 10674 11452
rect 10610 11392 10674 11396
rect 10690 11452 10754 11456
rect 10690 11396 10694 11452
rect 10694 11396 10750 11452
rect 10750 11396 10754 11452
rect 10690 11392 10754 11396
rect 10770 11452 10834 11456
rect 10770 11396 10774 11452
rect 10774 11396 10830 11452
rect 10830 11396 10834 11452
rect 10770 11392 10834 11396
rect 10850 11452 10914 11456
rect 10850 11396 10854 11452
rect 10854 11396 10910 11452
rect 10910 11396 10914 11452
rect 10850 11392 10914 11396
rect 17049 11452 17113 11456
rect 17049 11396 17053 11452
rect 17053 11396 17109 11452
rect 17109 11396 17113 11452
rect 17049 11392 17113 11396
rect 17129 11452 17193 11456
rect 17129 11396 17133 11452
rect 17133 11396 17189 11452
rect 17189 11396 17193 11452
rect 17129 11392 17193 11396
rect 17209 11452 17273 11456
rect 17209 11396 17213 11452
rect 17213 11396 17269 11452
rect 17269 11396 17273 11452
rect 17209 11392 17273 11396
rect 17289 11452 17353 11456
rect 17289 11396 17293 11452
rect 17293 11396 17349 11452
rect 17349 11396 17353 11452
rect 17289 11392 17353 11396
rect 23488 11452 23552 11456
rect 23488 11396 23492 11452
rect 23492 11396 23548 11452
rect 23548 11396 23552 11452
rect 23488 11392 23552 11396
rect 23568 11452 23632 11456
rect 23568 11396 23572 11452
rect 23572 11396 23628 11452
rect 23628 11396 23632 11452
rect 23568 11392 23632 11396
rect 23648 11452 23712 11456
rect 23648 11396 23652 11452
rect 23652 11396 23708 11452
rect 23708 11396 23712 11452
rect 23648 11392 23712 11396
rect 23728 11452 23792 11456
rect 23728 11396 23732 11452
rect 23732 11396 23788 11452
rect 23788 11396 23792 11452
rect 23728 11392 23792 11396
rect 4831 10908 4895 10912
rect 4831 10852 4835 10908
rect 4835 10852 4891 10908
rect 4891 10852 4895 10908
rect 4831 10848 4895 10852
rect 4911 10908 4975 10912
rect 4911 10852 4915 10908
rect 4915 10852 4971 10908
rect 4971 10852 4975 10908
rect 4911 10848 4975 10852
rect 4991 10908 5055 10912
rect 4991 10852 4995 10908
rect 4995 10852 5051 10908
rect 5051 10852 5055 10908
rect 4991 10848 5055 10852
rect 5071 10908 5135 10912
rect 5071 10852 5075 10908
rect 5075 10852 5131 10908
rect 5131 10852 5135 10908
rect 5071 10848 5135 10852
rect 11270 10908 11334 10912
rect 11270 10852 11274 10908
rect 11274 10852 11330 10908
rect 11330 10852 11334 10908
rect 11270 10848 11334 10852
rect 11350 10908 11414 10912
rect 11350 10852 11354 10908
rect 11354 10852 11410 10908
rect 11410 10852 11414 10908
rect 11350 10848 11414 10852
rect 11430 10908 11494 10912
rect 11430 10852 11434 10908
rect 11434 10852 11490 10908
rect 11490 10852 11494 10908
rect 11430 10848 11494 10852
rect 11510 10908 11574 10912
rect 11510 10852 11514 10908
rect 11514 10852 11570 10908
rect 11570 10852 11574 10908
rect 11510 10848 11574 10852
rect 17709 10908 17773 10912
rect 17709 10852 17713 10908
rect 17713 10852 17769 10908
rect 17769 10852 17773 10908
rect 17709 10848 17773 10852
rect 17789 10908 17853 10912
rect 17789 10852 17793 10908
rect 17793 10852 17849 10908
rect 17849 10852 17853 10908
rect 17789 10848 17853 10852
rect 17869 10908 17933 10912
rect 17869 10852 17873 10908
rect 17873 10852 17929 10908
rect 17929 10852 17933 10908
rect 17869 10848 17933 10852
rect 17949 10908 18013 10912
rect 17949 10852 17953 10908
rect 17953 10852 18009 10908
rect 18009 10852 18013 10908
rect 17949 10848 18013 10852
rect 24148 10908 24212 10912
rect 24148 10852 24152 10908
rect 24152 10852 24208 10908
rect 24208 10852 24212 10908
rect 24148 10848 24212 10852
rect 24228 10908 24292 10912
rect 24228 10852 24232 10908
rect 24232 10852 24288 10908
rect 24288 10852 24292 10908
rect 24228 10848 24292 10852
rect 24308 10908 24372 10912
rect 24308 10852 24312 10908
rect 24312 10852 24368 10908
rect 24368 10852 24372 10908
rect 24308 10848 24372 10852
rect 24388 10908 24452 10912
rect 24388 10852 24392 10908
rect 24392 10852 24448 10908
rect 24448 10852 24452 10908
rect 24388 10848 24452 10852
rect 4171 10364 4235 10368
rect 4171 10308 4175 10364
rect 4175 10308 4231 10364
rect 4231 10308 4235 10364
rect 4171 10304 4235 10308
rect 4251 10364 4315 10368
rect 4251 10308 4255 10364
rect 4255 10308 4311 10364
rect 4311 10308 4315 10364
rect 4251 10304 4315 10308
rect 4331 10364 4395 10368
rect 4331 10308 4335 10364
rect 4335 10308 4391 10364
rect 4391 10308 4395 10364
rect 4331 10304 4395 10308
rect 4411 10364 4475 10368
rect 4411 10308 4415 10364
rect 4415 10308 4471 10364
rect 4471 10308 4475 10364
rect 4411 10304 4475 10308
rect 10610 10364 10674 10368
rect 10610 10308 10614 10364
rect 10614 10308 10670 10364
rect 10670 10308 10674 10364
rect 10610 10304 10674 10308
rect 10690 10364 10754 10368
rect 10690 10308 10694 10364
rect 10694 10308 10750 10364
rect 10750 10308 10754 10364
rect 10690 10304 10754 10308
rect 10770 10364 10834 10368
rect 10770 10308 10774 10364
rect 10774 10308 10830 10364
rect 10830 10308 10834 10364
rect 10770 10304 10834 10308
rect 10850 10364 10914 10368
rect 10850 10308 10854 10364
rect 10854 10308 10910 10364
rect 10910 10308 10914 10364
rect 10850 10304 10914 10308
rect 17049 10364 17113 10368
rect 17049 10308 17053 10364
rect 17053 10308 17109 10364
rect 17109 10308 17113 10364
rect 17049 10304 17113 10308
rect 17129 10364 17193 10368
rect 17129 10308 17133 10364
rect 17133 10308 17189 10364
rect 17189 10308 17193 10364
rect 17129 10304 17193 10308
rect 17209 10364 17273 10368
rect 17209 10308 17213 10364
rect 17213 10308 17269 10364
rect 17269 10308 17273 10364
rect 17209 10304 17273 10308
rect 17289 10364 17353 10368
rect 17289 10308 17293 10364
rect 17293 10308 17349 10364
rect 17349 10308 17353 10364
rect 17289 10304 17353 10308
rect 23488 10364 23552 10368
rect 23488 10308 23492 10364
rect 23492 10308 23548 10364
rect 23548 10308 23552 10364
rect 23488 10304 23552 10308
rect 23568 10364 23632 10368
rect 23568 10308 23572 10364
rect 23572 10308 23628 10364
rect 23628 10308 23632 10364
rect 23568 10304 23632 10308
rect 23648 10364 23712 10368
rect 23648 10308 23652 10364
rect 23652 10308 23708 10364
rect 23708 10308 23712 10364
rect 23648 10304 23712 10308
rect 23728 10364 23792 10368
rect 23728 10308 23732 10364
rect 23732 10308 23788 10364
rect 23788 10308 23792 10364
rect 23728 10304 23792 10308
rect 4831 9820 4895 9824
rect 4831 9764 4835 9820
rect 4835 9764 4891 9820
rect 4891 9764 4895 9820
rect 4831 9760 4895 9764
rect 4911 9820 4975 9824
rect 4911 9764 4915 9820
rect 4915 9764 4971 9820
rect 4971 9764 4975 9820
rect 4911 9760 4975 9764
rect 4991 9820 5055 9824
rect 4991 9764 4995 9820
rect 4995 9764 5051 9820
rect 5051 9764 5055 9820
rect 4991 9760 5055 9764
rect 5071 9820 5135 9824
rect 5071 9764 5075 9820
rect 5075 9764 5131 9820
rect 5131 9764 5135 9820
rect 5071 9760 5135 9764
rect 11270 9820 11334 9824
rect 11270 9764 11274 9820
rect 11274 9764 11330 9820
rect 11330 9764 11334 9820
rect 11270 9760 11334 9764
rect 11350 9820 11414 9824
rect 11350 9764 11354 9820
rect 11354 9764 11410 9820
rect 11410 9764 11414 9820
rect 11350 9760 11414 9764
rect 11430 9820 11494 9824
rect 11430 9764 11434 9820
rect 11434 9764 11490 9820
rect 11490 9764 11494 9820
rect 11430 9760 11494 9764
rect 11510 9820 11574 9824
rect 11510 9764 11514 9820
rect 11514 9764 11570 9820
rect 11570 9764 11574 9820
rect 11510 9760 11574 9764
rect 17709 9820 17773 9824
rect 17709 9764 17713 9820
rect 17713 9764 17769 9820
rect 17769 9764 17773 9820
rect 17709 9760 17773 9764
rect 17789 9820 17853 9824
rect 17789 9764 17793 9820
rect 17793 9764 17849 9820
rect 17849 9764 17853 9820
rect 17789 9760 17853 9764
rect 17869 9820 17933 9824
rect 17869 9764 17873 9820
rect 17873 9764 17929 9820
rect 17929 9764 17933 9820
rect 17869 9760 17933 9764
rect 17949 9820 18013 9824
rect 17949 9764 17953 9820
rect 17953 9764 18009 9820
rect 18009 9764 18013 9820
rect 17949 9760 18013 9764
rect 24148 9820 24212 9824
rect 24148 9764 24152 9820
rect 24152 9764 24208 9820
rect 24208 9764 24212 9820
rect 24148 9760 24212 9764
rect 24228 9820 24292 9824
rect 24228 9764 24232 9820
rect 24232 9764 24288 9820
rect 24288 9764 24292 9820
rect 24228 9760 24292 9764
rect 24308 9820 24372 9824
rect 24308 9764 24312 9820
rect 24312 9764 24368 9820
rect 24368 9764 24372 9820
rect 24308 9760 24372 9764
rect 24388 9820 24452 9824
rect 24388 9764 24392 9820
rect 24392 9764 24448 9820
rect 24448 9764 24452 9820
rect 24388 9760 24452 9764
rect 4171 9276 4235 9280
rect 4171 9220 4175 9276
rect 4175 9220 4231 9276
rect 4231 9220 4235 9276
rect 4171 9216 4235 9220
rect 4251 9276 4315 9280
rect 4251 9220 4255 9276
rect 4255 9220 4311 9276
rect 4311 9220 4315 9276
rect 4251 9216 4315 9220
rect 4331 9276 4395 9280
rect 4331 9220 4335 9276
rect 4335 9220 4391 9276
rect 4391 9220 4395 9276
rect 4331 9216 4395 9220
rect 4411 9276 4475 9280
rect 4411 9220 4415 9276
rect 4415 9220 4471 9276
rect 4471 9220 4475 9276
rect 4411 9216 4475 9220
rect 10610 9276 10674 9280
rect 10610 9220 10614 9276
rect 10614 9220 10670 9276
rect 10670 9220 10674 9276
rect 10610 9216 10674 9220
rect 10690 9276 10754 9280
rect 10690 9220 10694 9276
rect 10694 9220 10750 9276
rect 10750 9220 10754 9276
rect 10690 9216 10754 9220
rect 10770 9276 10834 9280
rect 10770 9220 10774 9276
rect 10774 9220 10830 9276
rect 10830 9220 10834 9276
rect 10770 9216 10834 9220
rect 10850 9276 10914 9280
rect 10850 9220 10854 9276
rect 10854 9220 10910 9276
rect 10910 9220 10914 9276
rect 10850 9216 10914 9220
rect 17049 9276 17113 9280
rect 17049 9220 17053 9276
rect 17053 9220 17109 9276
rect 17109 9220 17113 9276
rect 17049 9216 17113 9220
rect 17129 9276 17193 9280
rect 17129 9220 17133 9276
rect 17133 9220 17189 9276
rect 17189 9220 17193 9276
rect 17129 9216 17193 9220
rect 17209 9276 17273 9280
rect 17209 9220 17213 9276
rect 17213 9220 17269 9276
rect 17269 9220 17273 9276
rect 17209 9216 17273 9220
rect 17289 9276 17353 9280
rect 17289 9220 17293 9276
rect 17293 9220 17349 9276
rect 17349 9220 17353 9276
rect 17289 9216 17353 9220
rect 23488 9276 23552 9280
rect 23488 9220 23492 9276
rect 23492 9220 23548 9276
rect 23548 9220 23552 9276
rect 23488 9216 23552 9220
rect 23568 9276 23632 9280
rect 23568 9220 23572 9276
rect 23572 9220 23628 9276
rect 23628 9220 23632 9276
rect 23568 9216 23632 9220
rect 23648 9276 23712 9280
rect 23648 9220 23652 9276
rect 23652 9220 23708 9276
rect 23708 9220 23712 9276
rect 23648 9216 23712 9220
rect 23728 9276 23792 9280
rect 23728 9220 23732 9276
rect 23732 9220 23788 9276
rect 23788 9220 23792 9276
rect 23728 9216 23792 9220
rect 4831 8732 4895 8736
rect 4831 8676 4835 8732
rect 4835 8676 4891 8732
rect 4891 8676 4895 8732
rect 4831 8672 4895 8676
rect 4911 8732 4975 8736
rect 4911 8676 4915 8732
rect 4915 8676 4971 8732
rect 4971 8676 4975 8732
rect 4911 8672 4975 8676
rect 4991 8732 5055 8736
rect 4991 8676 4995 8732
rect 4995 8676 5051 8732
rect 5051 8676 5055 8732
rect 4991 8672 5055 8676
rect 5071 8732 5135 8736
rect 5071 8676 5075 8732
rect 5075 8676 5131 8732
rect 5131 8676 5135 8732
rect 5071 8672 5135 8676
rect 11270 8732 11334 8736
rect 11270 8676 11274 8732
rect 11274 8676 11330 8732
rect 11330 8676 11334 8732
rect 11270 8672 11334 8676
rect 11350 8732 11414 8736
rect 11350 8676 11354 8732
rect 11354 8676 11410 8732
rect 11410 8676 11414 8732
rect 11350 8672 11414 8676
rect 11430 8732 11494 8736
rect 11430 8676 11434 8732
rect 11434 8676 11490 8732
rect 11490 8676 11494 8732
rect 11430 8672 11494 8676
rect 11510 8732 11574 8736
rect 11510 8676 11514 8732
rect 11514 8676 11570 8732
rect 11570 8676 11574 8732
rect 11510 8672 11574 8676
rect 17709 8732 17773 8736
rect 17709 8676 17713 8732
rect 17713 8676 17769 8732
rect 17769 8676 17773 8732
rect 17709 8672 17773 8676
rect 17789 8732 17853 8736
rect 17789 8676 17793 8732
rect 17793 8676 17849 8732
rect 17849 8676 17853 8732
rect 17789 8672 17853 8676
rect 17869 8732 17933 8736
rect 17869 8676 17873 8732
rect 17873 8676 17929 8732
rect 17929 8676 17933 8732
rect 17869 8672 17933 8676
rect 17949 8732 18013 8736
rect 17949 8676 17953 8732
rect 17953 8676 18009 8732
rect 18009 8676 18013 8732
rect 17949 8672 18013 8676
rect 24148 8732 24212 8736
rect 24148 8676 24152 8732
rect 24152 8676 24208 8732
rect 24208 8676 24212 8732
rect 24148 8672 24212 8676
rect 24228 8732 24292 8736
rect 24228 8676 24232 8732
rect 24232 8676 24288 8732
rect 24288 8676 24292 8732
rect 24228 8672 24292 8676
rect 24308 8732 24372 8736
rect 24308 8676 24312 8732
rect 24312 8676 24368 8732
rect 24368 8676 24372 8732
rect 24308 8672 24372 8676
rect 24388 8732 24452 8736
rect 24388 8676 24392 8732
rect 24392 8676 24448 8732
rect 24448 8676 24452 8732
rect 24388 8672 24452 8676
rect 4171 8188 4235 8192
rect 4171 8132 4175 8188
rect 4175 8132 4231 8188
rect 4231 8132 4235 8188
rect 4171 8128 4235 8132
rect 4251 8188 4315 8192
rect 4251 8132 4255 8188
rect 4255 8132 4311 8188
rect 4311 8132 4315 8188
rect 4251 8128 4315 8132
rect 4331 8188 4395 8192
rect 4331 8132 4335 8188
rect 4335 8132 4391 8188
rect 4391 8132 4395 8188
rect 4331 8128 4395 8132
rect 4411 8188 4475 8192
rect 4411 8132 4415 8188
rect 4415 8132 4471 8188
rect 4471 8132 4475 8188
rect 4411 8128 4475 8132
rect 10610 8188 10674 8192
rect 10610 8132 10614 8188
rect 10614 8132 10670 8188
rect 10670 8132 10674 8188
rect 10610 8128 10674 8132
rect 10690 8188 10754 8192
rect 10690 8132 10694 8188
rect 10694 8132 10750 8188
rect 10750 8132 10754 8188
rect 10690 8128 10754 8132
rect 10770 8188 10834 8192
rect 10770 8132 10774 8188
rect 10774 8132 10830 8188
rect 10830 8132 10834 8188
rect 10770 8128 10834 8132
rect 10850 8188 10914 8192
rect 10850 8132 10854 8188
rect 10854 8132 10910 8188
rect 10910 8132 10914 8188
rect 10850 8128 10914 8132
rect 17049 8188 17113 8192
rect 17049 8132 17053 8188
rect 17053 8132 17109 8188
rect 17109 8132 17113 8188
rect 17049 8128 17113 8132
rect 17129 8188 17193 8192
rect 17129 8132 17133 8188
rect 17133 8132 17189 8188
rect 17189 8132 17193 8188
rect 17129 8128 17193 8132
rect 17209 8188 17273 8192
rect 17209 8132 17213 8188
rect 17213 8132 17269 8188
rect 17269 8132 17273 8188
rect 17209 8128 17273 8132
rect 17289 8188 17353 8192
rect 17289 8132 17293 8188
rect 17293 8132 17349 8188
rect 17349 8132 17353 8188
rect 17289 8128 17353 8132
rect 23488 8188 23552 8192
rect 23488 8132 23492 8188
rect 23492 8132 23548 8188
rect 23548 8132 23552 8188
rect 23488 8128 23552 8132
rect 23568 8188 23632 8192
rect 23568 8132 23572 8188
rect 23572 8132 23628 8188
rect 23628 8132 23632 8188
rect 23568 8128 23632 8132
rect 23648 8188 23712 8192
rect 23648 8132 23652 8188
rect 23652 8132 23708 8188
rect 23708 8132 23712 8188
rect 23648 8128 23712 8132
rect 23728 8188 23792 8192
rect 23728 8132 23732 8188
rect 23732 8132 23788 8188
rect 23788 8132 23792 8188
rect 23728 8128 23792 8132
rect 4831 7644 4895 7648
rect 4831 7588 4835 7644
rect 4835 7588 4891 7644
rect 4891 7588 4895 7644
rect 4831 7584 4895 7588
rect 4911 7644 4975 7648
rect 4911 7588 4915 7644
rect 4915 7588 4971 7644
rect 4971 7588 4975 7644
rect 4911 7584 4975 7588
rect 4991 7644 5055 7648
rect 4991 7588 4995 7644
rect 4995 7588 5051 7644
rect 5051 7588 5055 7644
rect 4991 7584 5055 7588
rect 5071 7644 5135 7648
rect 5071 7588 5075 7644
rect 5075 7588 5131 7644
rect 5131 7588 5135 7644
rect 5071 7584 5135 7588
rect 11270 7644 11334 7648
rect 11270 7588 11274 7644
rect 11274 7588 11330 7644
rect 11330 7588 11334 7644
rect 11270 7584 11334 7588
rect 11350 7644 11414 7648
rect 11350 7588 11354 7644
rect 11354 7588 11410 7644
rect 11410 7588 11414 7644
rect 11350 7584 11414 7588
rect 11430 7644 11494 7648
rect 11430 7588 11434 7644
rect 11434 7588 11490 7644
rect 11490 7588 11494 7644
rect 11430 7584 11494 7588
rect 11510 7644 11574 7648
rect 11510 7588 11514 7644
rect 11514 7588 11570 7644
rect 11570 7588 11574 7644
rect 11510 7584 11574 7588
rect 17709 7644 17773 7648
rect 17709 7588 17713 7644
rect 17713 7588 17769 7644
rect 17769 7588 17773 7644
rect 17709 7584 17773 7588
rect 17789 7644 17853 7648
rect 17789 7588 17793 7644
rect 17793 7588 17849 7644
rect 17849 7588 17853 7644
rect 17789 7584 17853 7588
rect 17869 7644 17933 7648
rect 17869 7588 17873 7644
rect 17873 7588 17929 7644
rect 17929 7588 17933 7644
rect 17869 7584 17933 7588
rect 17949 7644 18013 7648
rect 17949 7588 17953 7644
rect 17953 7588 18009 7644
rect 18009 7588 18013 7644
rect 17949 7584 18013 7588
rect 24148 7644 24212 7648
rect 24148 7588 24152 7644
rect 24152 7588 24208 7644
rect 24208 7588 24212 7644
rect 24148 7584 24212 7588
rect 24228 7644 24292 7648
rect 24228 7588 24232 7644
rect 24232 7588 24288 7644
rect 24288 7588 24292 7644
rect 24228 7584 24292 7588
rect 24308 7644 24372 7648
rect 24308 7588 24312 7644
rect 24312 7588 24368 7644
rect 24368 7588 24372 7644
rect 24308 7584 24372 7588
rect 24388 7644 24452 7648
rect 24388 7588 24392 7644
rect 24392 7588 24448 7644
rect 24448 7588 24452 7644
rect 24388 7584 24452 7588
rect 4171 7100 4235 7104
rect 4171 7044 4175 7100
rect 4175 7044 4231 7100
rect 4231 7044 4235 7100
rect 4171 7040 4235 7044
rect 4251 7100 4315 7104
rect 4251 7044 4255 7100
rect 4255 7044 4311 7100
rect 4311 7044 4315 7100
rect 4251 7040 4315 7044
rect 4331 7100 4395 7104
rect 4331 7044 4335 7100
rect 4335 7044 4391 7100
rect 4391 7044 4395 7100
rect 4331 7040 4395 7044
rect 4411 7100 4475 7104
rect 4411 7044 4415 7100
rect 4415 7044 4471 7100
rect 4471 7044 4475 7100
rect 4411 7040 4475 7044
rect 10610 7100 10674 7104
rect 10610 7044 10614 7100
rect 10614 7044 10670 7100
rect 10670 7044 10674 7100
rect 10610 7040 10674 7044
rect 10690 7100 10754 7104
rect 10690 7044 10694 7100
rect 10694 7044 10750 7100
rect 10750 7044 10754 7100
rect 10690 7040 10754 7044
rect 10770 7100 10834 7104
rect 10770 7044 10774 7100
rect 10774 7044 10830 7100
rect 10830 7044 10834 7100
rect 10770 7040 10834 7044
rect 10850 7100 10914 7104
rect 10850 7044 10854 7100
rect 10854 7044 10910 7100
rect 10910 7044 10914 7100
rect 10850 7040 10914 7044
rect 17049 7100 17113 7104
rect 17049 7044 17053 7100
rect 17053 7044 17109 7100
rect 17109 7044 17113 7100
rect 17049 7040 17113 7044
rect 17129 7100 17193 7104
rect 17129 7044 17133 7100
rect 17133 7044 17189 7100
rect 17189 7044 17193 7100
rect 17129 7040 17193 7044
rect 17209 7100 17273 7104
rect 17209 7044 17213 7100
rect 17213 7044 17269 7100
rect 17269 7044 17273 7100
rect 17209 7040 17273 7044
rect 17289 7100 17353 7104
rect 17289 7044 17293 7100
rect 17293 7044 17349 7100
rect 17349 7044 17353 7100
rect 17289 7040 17353 7044
rect 23488 7100 23552 7104
rect 23488 7044 23492 7100
rect 23492 7044 23548 7100
rect 23548 7044 23552 7100
rect 23488 7040 23552 7044
rect 23568 7100 23632 7104
rect 23568 7044 23572 7100
rect 23572 7044 23628 7100
rect 23628 7044 23632 7100
rect 23568 7040 23632 7044
rect 23648 7100 23712 7104
rect 23648 7044 23652 7100
rect 23652 7044 23708 7100
rect 23708 7044 23712 7100
rect 23648 7040 23712 7044
rect 23728 7100 23792 7104
rect 23728 7044 23732 7100
rect 23732 7044 23788 7100
rect 23788 7044 23792 7100
rect 23728 7040 23792 7044
rect 4831 6556 4895 6560
rect 4831 6500 4835 6556
rect 4835 6500 4891 6556
rect 4891 6500 4895 6556
rect 4831 6496 4895 6500
rect 4911 6556 4975 6560
rect 4911 6500 4915 6556
rect 4915 6500 4971 6556
rect 4971 6500 4975 6556
rect 4911 6496 4975 6500
rect 4991 6556 5055 6560
rect 4991 6500 4995 6556
rect 4995 6500 5051 6556
rect 5051 6500 5055 6556
rect 4991 6496 5055 6500
rect 5071 6556 5135 6560
rect 5071 6500 5075 6556
rect 5075 6500 5131 6556
rect 5131 6500 5135 6556
rect 5071 6496 5135 6500
rect 11270 6556 11334 6560
rect 11270 6500 11274 6556
rect 11274 6500 11330 6556
rect 11330 6500 11334 6556
rect 11270 6496 11334 6500
rect 11350 6556 11414 6560
rect 11350 6500 11354 6556
rect 11354 6500 11410 6556
rect 11410 6500 11414 6556
rect 11350 6496 11414 6500
rect 11430 6556 11494 6560
rect 11430 6500 11434 6556
rect 11434 6500 11490 6556
rect 11490 6500 11494 6556
rect 11430 6496 11494 6500
rect 11510 6556 11574 6560
rect 11510 6500 11514 6556
rect 11514 6500 11570 6556
rect 11570 6500 11574 6556
rect 11510 6496 11574 6500
rect 17709 6556 17773 6560
rect 17709 6500 17713 6556
rect 17713 6500 17769 6556
rect 17769 6500 17773 6556
rect 17709 6496 17773 6500
rect 17789 6556 17853 6560
rect 17789 6500 17793 6556
rect 17793 6500 17849 6556
rect 17849 6500 17853 6556
rect 17789 6496 17853 6500
rect 17869 6556 17933 6560
rect 17869 6500 17873 6556
rect 17873 6500 17929 6556
rect 17929 6500 17933 6556
rect 17869 6496 17933 6500
rect 17949 6556 18013 6560
rect 17949 6500 17953 6556
rect 17953 6500 18009 6556
rect 18009 6500 18013 6556
rect 17949 6496 18013 6500
rect 24148 6556 24212 6560
rect 24148 6500 24152 6556
rect 24152 6500 24208 6556
rect 24208 6500 24212 6556
rect 24148 6496 24212 6500
rect 24228 6556 24292 6560
rect 24228 6500 24232 6556
rect 24232 6500 24288 6556
rect 24288 6500 24292 6556
rect 24228 6496 24292 6500
rect 24308 6556 24372 6560
rect 24308 6500 24312 6556
rect 24312 6500 24368 6556
rect 24368 6500 24372 6556
rect 24308 6496 24372 6500
rect 24388 6556 24452 6560
rect 24388 6500 24392 6556
rect 24392 6500 24448 6556
rect 24448 6500 24452 6556
rect 24388 6496 24452 6500
rect 4171 6012 4235 6016
rect 4171 5956 4175 6012
rect 4175 5956 4231 6012
rect 4231 5956 4235 6012
rect 4171 5952 4235 5956
rect 4251 6012 4315 6016
rect 4251 5956 4255 6012
rect 4255 5956 4311 6012
rect 4311 5956 4315 6012
rect 4251 5952 4315 5956
rect 4331 6012 4395 6016
rect 4331 5956 4335 6012
rect 4335 5956 4391 6012
rect 4391 5956 4395 6012
rect 4331 5952 4395 5956
rect 4411 6012 4475 6016
rect 4411 5956 4415 6012
rect 4415 5956 4471 6012
rect 4471 5956 4475 6012
rect 4411 5952 4475 5956
rect 10610 6012 10674 6016
rect 10610 5956 10614 6012
rect 10614 5956 10670 6012
rect 10670 5956 10674 6012
rect 10610 5952 10674 5956
rect 10690 6012 10754 6016
rect 10690 5956 10694 6012
rect 10694 5956 10750 6012
rect 10750 5956 10754 6012
rect 10690 5952 10754 5956
rect 10770 6012 10834 6016
rect 10770 5956 10774 6012
rect 10774 5956 10830 6012
rect 10830 5956 10834 6012
rect 10770 5952 10834 5956
rect 10850 6012 10914 6016
rect 10850 5956 10854 6012
rect 10854 5956 10910 6012
rect 10910 5956 10914 6012
rect 10850 5952 10914 5956
rect 17049 6012 17113 6016
rect 17049 5956 17053 6012
rect 17053 5956 17109 6012
rect 17109 5956 17113 6012
rect 17049 5952 17113 5956
rect 17129 6012 17193 6016
rect 17129 5956 17133 6012
rect 17133 5956 17189 6012
rect 17189 5956 17193 6012
rect 17129 5952 17193 5956
rect 17209 6012 17273 6016
rect 17209 5956 17213 6012
rect 17213 5956 17269 6012
rect 17269 5956 17273 6012
rect 17209 5952 17273 5956
rect 17289 6012 17353 6016
rect 17289 5956 17293 6012
rect 17293 5956 17349 6012
rect 17349 5956 17353 6012
rect 17289 5952 17353 5956
rect 23488 6012 23552 6016
rect 23488 5956 23492 6012
rect 23492 5956 23548 6012
rect 23548 5956 23552 6012
rect 23488 5952 23552 5956
rect 23568 6012 23632 6016
rect 23568 5956 23572 6012
rect 23572 5956 23628 6012
rect 23628 5956 23632 6012
rect 23568 5952 23632 5956
rect 23648 6012 23712 6016
rect 23648 5956 23652 6012
rect 23652 5956 23708 6012
rect 23708 5956 23712 6012
rect 23648 5952 23712 5956
rect 23728 6012 23792 6016
rect 23728 5956 23732 6012
rect 23732 5956 23788 6012
rect 23788 5956 23792 6012
rect 23728 5952 23792 5956
rect 4831 5468 4895 5472
rect 4831 5412 4835 5468
rect 4835 5412 4891 5468
rect 4891 5412 4895 5468
rect 4831 5408 4895 5412
rect 4911 5468 4975 5472
rect 4911 5412 4915 5468
rect 4915 5412 4971 5468
rect 4971 5412 4975 5468
rect 4911 5408 4975 5412
rect 4991 5468 5055 5472
rect 4991 5412 4995 5468
rect 4995 5412 5051 5468
rect 5051 5412 5055 5468
rect 4991 5408 5055 5412
rect 5071 5468 5135 5472
rect 5071 5412 5075 5468
rect 5075 5412 5131 5468
rect 5131 5412 5135 5468
rect 5071 5408 5135 5412
rect 11270 5468 11334 5472
rect 11270 5412 11274 5468
rect 11274 5412 11330 5468
rect 11330 5412 11334 5468
rect 11270 5408 11334 5412
rect 11350 5468 11414 5472
rect 11350 5412 11354 5468
rect 11354 5412 11410 5468
rect 11410 5412 11414 5468
rect 11350 5408 11414 5412
rect 11430 5468 11494 5472
rect 11430 5412 11434 5468
rect 11434 5412 11490 5468
rect 11490 5412 11494 5468
rect 11430 5408 11494 5412
rect 11510 5468 11574 5472
rect 11510 5412 11514 5468
rect 11514 5412 11570 5468
rect 11570 5412 11574 5468
rect 11510 5408 11574 5412
rect 17709 5468 17773 5472
rect 17709 5412 17713 5468
rect 17713 5412 17769 5468
rect 17769 5412 17773 5468
rect 17709 5408 17773 5412
rect 17789 5468 17853 5472
rect 17789 5412 17793 5468
rect 17793 5412 17849 5468
rect 17849 5412 17853 5468
rect 17789 5408 17853 5412
rect 17869 5468 17933 5472
rect 17869 5412 17873 5468
rect 17873 5412 17929 5468
rect 17929 5412 17933 5468
rect 17869 5408 17933 5412
rect 17949 5468 18013 5472
rect 17949 5412 17953 5468
rect 17953 5412 18009 5468
rect 18009 5412 18013 5468
rect 17949 5408 18013 5412
rect 24148 5468 24212 5472
rect 24148 5412 24152 5468
rect 24152 5412 24208 5468
rect 24208 5412 24212 5468
rect 24148 5408 24212 5412
rect 24228 5468 24292 5472
rect 24228 5412 24232 5468
rect 24232 5412 24288 5468
rect 24288 5412 24292 5468
rect 24228 5408 24292 5412
rect 24308 5468 24372 5472
rect 24308 5412 24312 5468
rect 24312 5412 24368 5468
rect 24368 5412 24372 5468
rect 24308 5408 24372 5412
rect 24388 5468 24452 5472
rect 24388 5412 24392 5468
rect 24392 5412 24448 5468
rect 24448 5412 24452 5468
rect 24388 5408 24452 5412
rect 4171 4924 4235 4928
rect 4171 4868 4175 4924
rect 4175 4868 4231 4924
rect 4231 4868 4235 4924
rect 4171 4864 4235 4868
rect 4251 4924 4315 4928
rect 4251 4868 4255 4924
rect 4255 4868 4311 4924
rect 4311 4868 4315 4924
rect 4251 4864 4315 4868
rect 4331 4924 4395 4928
rect 4331 4868 4335 4924
rect 4335 4868 4391 4924
rect 4391 4868 4395 4924
rect 4331 4864 4395 4868
rect 4411 4924 4475 4928
rect 4411 4868 4415 4924
rect 4415 4868 4471 4924
rect 4471 4868 4475 4924
rect 4411 4864 4475 4868
rect 10610 4924 10674 4928
rect 10610 4868 10614 4924
rect 10614 4868 10670 4924
rect 10670 4868 10674 4924
rect 10610 4864 10674 4868
rect 10690 4924 10754 4928
rect 10690 4868 10694 4924
rect 10694 4868 10750 4924
rect 10750 4868 10754 4924
rect 10690 4864 10754 4868
rect 10770 4924 10834 4928
rect 10770 4868 10774 4924
rect 10774 4868 10830 4924
rect 10830 4868 10834 4924
rect 10770 4864 10834 4868
rect 10850 4924 10914 4928
rect 10850 4868 10854 4924
rect 10854 4868 10910 4924
rect 10910 4868 10914 4924
rect 10850 4864 10914 4868
rect 17049 4924 17113 4928
rect 17049 4868 17053 4924
rect 17053 4868 17109 4924
rect 17109 4868 17113 4924
rect 17049 4864 17113 4868
rect 17129 4924 17193 4928
rect 17129 4868 17133 4924
rect 17133 4868 17189 4924
rect 17189 4868 17193 4924
rect 17129 4864 17193 4868
rect 17209 4924 17273 4928
rect 17209 4868 17213 4924
rect 17213 4868 17269 4924
rect 17269 4868 17273 4924
rect 17209 4864 17273 4868
rect 17289 4924 17353 4928
rect 17289 4868 17293 4924
rect 17293 4868 17349 4924
rect 17349 4868 17353 4924
rect 17289 4864 17353 4868
rect 23488 4924 23552 4928
rect 23488 4868 23492 4924
rect 23492 4868 23548 4924
rect 23548 4868 23552 4924
rect 23488 4864 23552 4868
rect 23568 4924 23632 4928
rect 23568 4868 23572 4924
rect 23572 4868 23628 4924
rect 23628 4868 23632 4924
rect 23568 4864 23632 4868
rect 23648 4924 23712 4928
rect 23648 4868 23652 4924
rect 23652 4868 23708 4924
rect 23708 4868 23712 4924
rect 23648 4864 23712 4868
rect 23728 4924 23792 4928
rect 23728 4868 23732 4924
rect 23732 4868 23788 4924
rect 23788 4868 23792 4924
rect 23728 4864 23792 4868
rect 4831 4380 4895 4384
rect 4831 4324 4835 4380
rect 4835 4324 4891 4380
rect 4891 4324 4895 4380
rect 4831 4320 4895 4324
rect 4911 4380 4975 4384
rect 4911 4324 4915 4380
rect 4915 4324 4971 4380
rect 4971 4324 4975 4380
rect 4911 4320 4975 4324
rect 4991 4380 5055 4384
rect 4991 4324 4995 4380
rect 4995 4324 5051 4380
rect 5051 4324 5055 4380
rect 4991 4320 5055 4324
rect 5071 4380 5135 4384
rect 5071 4324 5075 4380
rect 5075 4324 5131 4380
rect 5131 4324 5135 4380
rect 5071 4320 5135 4324
rect 11270 4380 11334 4384
rect 11270 4324 11274 4380
rect 11274 4324 11330 4380
rect 11330 4324 11334 4380
rect 11270 4320 11334 4324
rect 11350 4380 11414 4384
rect 11350 4324 11354 4380
rect 11354 4324 11410 4380
rect 11410 4324 11414 4380
rect 11350 4320 11414 4324
rect 11430 4380 11494 4384
rect 11430 4324 11434 4380
rect 11434 4324 11490 4380
rect 11490 4324 11494 4380
rect 11430 4320 11494 4324
rect 11510 4380 11574 4384
rect 11510 4324 11514 4380
rect 11514 4324 11570 4380
rect 11570 4324 11574 4380
rect 11510 4320 11574 4324
rect 17709 4380 17773 4384
rect 17709 4324 17713 4380
rect 17713 4324 17769 4380
rect 17769 4324 17773 4380
rect 17709 4320 17773 4324
rect 17789 4380 17853 4384
rect 17789 4324 17793 4380
rect 17793 4324 17849 4380
rect 17849 4324 17853 4380
rect 17789 4320 17853 4324
rect 17869 4380 17933 4384
rect 17869 4324 17873 4380
rect 17873 4324 17929 4380
rect 17929 4324 17933 4380
rect 17869 4320 17933 4324
rect 17949 4380 18013 4384
rect 17949 4324 17953 4380
rect 17953 4324 18009 4380
rect 18009 4324 18013 4380
rect 17949 4320 18013 4324
rect 24148 4380 24212 4384
rect 24148 4324 24152 4380
rect 24152 4324 24208 4380
rect 24208 4324 24212 4380
rect 24148 4320 24212 4324
rect 24228 4380 24292 4384
rect 24228 4324 24232 4380
rect 24232 4324 24288 4380
rect 24288 4324 24292 4380
rect 24228 4320 24292 4324
rect 24308 4380 24372 4384
rect 24308 4324 24312 4380
rect 24312 4324 24368 4380
rect 24368 4324 24372 4380
rect 24308 4320 24372 4324
rect 24388 4380 24452 4384
rect 24388 4324 24392 4380
rect 24392 4324 24448 4380
rect 24448 4324 24452 4380
rect 24388 4320 24452 4324
rect 4171 3836 4235 3840
rect 4171 3780 4175 3836
rect 4175 3780 4231 3836
rect 4231 3780 4235 3836
rect 4171 3776 4235 3780
rect 4251 3836 4315 3840
rect 4251 3780 4255 3836
rect 4255 3780 4311 3836
rect 4311 3780 4315 3836
rect 4251 3776 4315 3780
rect 4331 3836 4395 3840
rect 4331 3780 4335 3836
rect 4335 3780 4391 3836
rect 4391 3780 4395 3836
rect 4331 3776 4395 3780
rect 4411 3836 4475 3840
rect 4411 3780 4415 3836
rect 4415 3780 4471 3836
rect 4471 3780 4475 3836
rect 4411 3776 4475 3780
rect 10610 3836 10674 3840
rect 10610 3780 10614 3836
rect 10614 3780 10670 3836
rect 10670 3780 10674 3836
rect 10610 3776 10674 3780
rect 10690 3836 10754 3840
rect 10690 3780 10694 3836
rect 10694 3780 10750 3836
rect 10750 3780 10754 3836
rect 10690 3776 10754 3780
rect 10770 3836 10834 3840
rect 10770 3780 10774 3836
rect 10774 3780 10830 3836
rect 10830 3780 10834 3836
rect 10770 3776 10834 3780
rect 10850 3836 10914 3840
rect 10850 3780 10854 3836
rect 10854 3780 10910 3836
rect 10910 3780 10914 3836
rect 10850 3776 10914 3780
rect 17049 3836 17113 3840
rect 17049 3780 17053 3836
rect 17053 3780 17109 3836
rect 17109 3780 17113 3836
rect 17049 3776 17113 3780
rect 17129 3836 17193 3840
rect 17129 3780 17133 3836
rect 17133 3780 17189 3836
rect 17189 3780 17193 3836
rect 17129 3776 17193 3780
rect 17209 3836 17273 3840
rect 17209 3780 17213 3836
rect 17213 3780 17269 3836
rect 17269 3780 17273 3836
rect 17209 3776 17273 3780
rect 17289 3836 17353 3840
rect 17289 3780 17293 3836
rect 17293 3780 17349 3836
rect 17349 3780 17353 3836
rect 17289 3776 17353 3780
rect 23488 3836 23552 3840
rect 23488 3780 23492 3836
rect 23492 3780 23548 3836
rect 23548 3780 23552 3836
rect 23488 3776 23552 3780
rect 23568 3836 23632 3840
rect 23568 3780 23572 3836
rect 23572 3780 23628 3836
rect 23628 3780 23632 3836
rect 23568 3776 23632 3780
rect 23648 3836 23712 3840
rect 23648 3780 23652 3836
rect 23652 3780 23708 3836
rect 23708 3780 23712 3836
rect 23648 3776 23712 3780
rect 23728 3836 23792 3840
rect 23728 3780 23732 3836
rect 23732 3780 23788 3836
rect 23788 3780 23792 3836
rect 23728 3776 23792 3780
rect 4831 3292 4895 3296
rect 4831 3236 4835 3292
rect 4835 3236 4891 3292
rect 4891 3236 4895 3292
rect 4831 3232 4895 3236
rect 4911 3292 4975 3296
rect 4911 3236 4915 3292
rect 4915 3236 4971 3292
rect 4971 3236 4975 3292
rect 4911 3232 4975 3236
rect 4991 3292 5055 3296
rect 4991 3236 4995 3292
rect 4995 3236 5051 3292
rect 5051 3236 5055 3292
rect 4991 3232 5055 3236
rect 5071 3292 5135 3296
rect 5071 3236 5075 3292
rect 5075 3236 5131 3292
rect 5131 3236 5135 3292
rect 5071 3232 5135 3236
rect 11270 3292 11334 3296
rect 11270 3236 11274 3292
rect 11274 3236 11330 3292
rect 11330 3236 11334 3292
rect 11270 3232 11334 3236
rect 11350 3292 11414 3296
rect 11350 3236 11354 3292
rect 11354 3236 11410 3292
rect 11410 3236 11414 3292
rect 11350 3232 11414 3236
rect 11430 3292 11494 3296
rect 11430 3236 11434 3292
rect 11434 3236 11490 3292
rect 11490 3236 11494 3292
rect 11430 3232 11494 3236
rect 11510 3292 11574 3296
rect 11510 3236 11514 3292
rect 11514 3236 11570 3292
rect 11570 3236 11574 3292
rect 11510 3232 11574 3236
rect 17709 3292 17773 3296
rect 17709 3236 17713 3292
rect 17713 3236 17769 3292
rect 17769 3236 17773 3292
rect 17709 3232 17773 3236
rect 17789 3292 17853 3296
rect 17789 3236 17793 3292
rect 17793 3236 17849 3292
rect 17849 3236 17853 3292
rect 17789 3232 17853 3236
rect 17869 3292 17933 3296
rect 17869 3236 17873 3292
rect 17873 3236 17929 3292
rect 17929 3236 17933 3292
rect 17869 3232 17933 3236
rect 17949 3292 18013 3296
rect 17949 3236 17953 3292
rect 17953 3236 18009 3292
rect 18009 3236 18013 3292
rect 17949 3232 18013 3236
rect 24148 3292 24212 3296
rect 24148 3236 24152 3292
rect 24152 3236 24208 3292
rect 24208 3236 24212 3292
rect 24148 3232 24212 3236
rect 24228 3292 24292 3296
rect 24228 3236 24232 3292
rect 24232 3236 24288 3292
rect 24288 3236 24292 3292
rect 24228 3232 24292 3236
rect 24308 3292 24372 3296
rect 24308 3236 24312 3292
rect 24312 3236 24368 3292
rect 24368 3236 24372 3292
rect 24308 3232 24372 3236
rect 24388 3292 24452 3296
rect 24388 3236 24392 3292
rect 24392 3236 24448 3292
rect 24448 3236 24452 3292
rect 24388 3232 24452 3236
rect 4171 2748 4235 2752
rect 4171 2692 4175 2748
rect 4175 2692 4231 2748
rect 4231 2692 4235 2748
rect 4171 2688 4235 2692
rect 4251 2748 4315 2752
rect 4251 2692 4255 2748
rect 4255 2692 4311 2748
rect 4311 2692 4315 2748
rect 4251 2688 4315 2692
rect 4331 2748 4395 2752
rect 4331 2692 4335 2748
rect 4335 2692 4391 2748
rect 4391 2692 4395 2748
rect 4331 2688 4395 2692
rect 4411 2748 4475 2752
rect 4411 2692 4415 2748
rect 4415 2692 4471 2748
rect 4471 2692 4475 2748
rect 4411 2688 4475 2692
rect 10610 2748 10674 2752
rect 10610 2692 10614 2748
rect 10614 2692 10670 2748
rect 10670 2692 10674 2748
rect 10610 2688 10674 2692
rect 10690 2748 10754 2752
rect 10690 2692 10694 2748
rect 10694 2692 10750 2748
rect 10750 2692 10754 2748
rect 10690 2688 10754 2692
rect 10770 2748 10834 2752
rect 10770 2692 10774 2748
rect 10774 2692 10830 2748
rect 10830 2692 10834 2748
rect 10770 2688 10834 2692
rect 10850 2748 10914 2752
rect 10850 2692 10854 2748
rect 10854 2692 10910 2748
rect 10910 2692 10914 2748
rect 10850 2688 10914 2692
rect 17049 2748 17113 2752
rect 17049 2692 17053 2748
rect 17053 2692 17109 2748
rect 17109 2692 17113 2748
rect 17049 2688 17113 2692
rect 17129 2748 17193 2752
rect 17129 2692 17133 2748
rect 17133 2692 17189 2748
rect 17189 2692 17193 2748
rect 17129 2688 17193 2692
rect 17209 2748 17273 2752
rect 17209 2692 17213 2748
rect 17213 2692 17269 2748
rect 17269 2692 17273 2748
rect 17209 2688 17273 2692
rect 17289 2748 17353 2752
rect 17289 2692 17293 2748
rect 17293 2692 17349 2748
rect 17349 2692 17353 2748
rect 17289 2688 17353 2692
rect 23488 2748 23552 2752
rect 23488 2692 23492 2748
rect 23492 2692 23548 2748
rect 23548 2692 23552 2748
rect 23488 2688 23552 2692
rect 23568 2748 23632 2752
rect 23568 2692 23572 2748
rect 23572 2692 23628 2748
rect 23628 2692 23632 2748
rect 23568 2688 23632 2692
rect 23648 2748 23712 2752
rect 23648 2692 23652 2748
rect 23652 2692 23708 2748
rect 23708 2692 23712 2748
rect 23648 2688 23712 2692
rect 23728 2748 23792 2752
rect 23728 2692 23732 2748
rect 23732 2692 23788 2748
rect 23788 2692 23792 2748
rect 23728 2688 23792 2692
rect 4831 2204 4895 2208
rect 4831 2148 4835 2204
rect 4835 2148 4891 2204
rect 4891 2148 4895 2204
rect 4831 2144 4895 2148
rect 4911 2204 4975 2208
rect 4911 2148 4915 2204
rect 4915 2148 4971 2204
rect 4971 2148 4975 2204
rect 4911 2144 4975 2148
rect 4991 2204 5055 2208
rect 4991 2148 4995 2204
rect 4995 2148 5051 2204
rect 5051 2148 5055 2204
rect 4991 2144 5055 2148
rect 5071 2204 5135 2208
rect 5071 2148 5075 2204
rect 5075 2148 5131 2204
rect 5131 2148 5135 2204
rect 5071 2144 5135 2148
rect 11270 2204 11334 2208
rect 11270 2148 11274 2204
rect 11274 2148 11330 2204
rect 11330 2148 11334 2204
rect 11270 2144 11334 2148
rect 11350 2204 11414 2208
rect 11350 2148 11354 2204
rect 11354 2148 11410 2204
rect 11410 2148 11414 2204
rect 11350 2144 11414 2148
rect 11430 2204 11494 2208
rect 11430 2148 11434 2204
rect 11434 2148 11490 2204
rect 11490 2148 11494 2204
rect 11430 2144 11494 2148
rect 11510 2204 11574 2208
rect 11510 2148 11514 2204
rect 11514 2148 11570 2204
rect 11570 2148 11574 2204
rect 11510 2144 11574 2148
rect 17709 2204 17773 2208
rect 17709 2148 17713 2204
rect 17713 2148 17769 2204
rect 17769 2148 17773 2204
rect 17709 2144 17773 2148
rect 17789 2204 17853 2208
rect 17789 2148 17793 2204
rect 17793 2148 17849 2204
rect 17849 2148 17853 2204
rect 17789 2144 17853 2148
rect 17869 2204 17933 2208
rect 17869 2148 17873 2204
rect 17873 2148 17929 2204
rect 17929 2148 17933 2204
rect 17869 2144 17933 2148
rect 17949 2204 18013 2208
rect 17949 2148 17953 2204
rect 17953 2148 18009 2204
rect 18009 2148 18013 2204
rect 17949 2144 18013 2148
rect 24148 2204 24212 2208
rect 24148 2148 24152 2204
rect 24152 2148 24208 2204
rect 24208 2148 24212 2204
rect 24148 2144 24212 2148
rect 24228 2204 24292 2208
rect 24228 2148 24232 2204
rect 24232 2148 24288 2204
rect 24288 2148 24292 2204
rect 24228 2144 24292 2148
rect 24308 2204 24372 2208
rect 24308 2148 24312 2204
rect 24312 2148 24368 2204
rect 24368 2148 24372 2204
rect 24308 2144 24372 2148
rect 24388 2204 24452 2208
rect 24388 2148 24392 2204
rect 24392 2148 24448 2204
rect 24448 2148 24452 2204
rect 24388 2144 24452 2148
<< metal4 >>
rect 4163 27776 4483 27792
rect 4163 27712 4171 27776
rect 4235 27712 4251 27776
rect 4315 27712 4331 27776
rect 4395 27712 4411 27776
rect 4475 27712 4483 27776
rect 4163 26688 4483 27712
rect 4163 26624 4171 26688
rect 4235 26624 4251 26688
rect 4315 26624 4331 26688
rect 4395 26624 4411 26688
rect 4475 26624 4483 26688
rect 4163 25600 4483 26624
rect 4163 25536 4171 25600
rect 4235 25536 4251 25600
rect 4315 25536 4331 25600
rect 4395 25536 4411 25600
rect 4475 25536 4483 25600
rect 4163 24666 4483 25536
rect 4163 24512 4205 24666
rect 4441 24512 4483 24666
rect 4163 24448 4171 24512
rect 4475 24448 4483 24512
rect 4163 24430 4205 24448
rect 4441 24430 4483 24448
rect 4163 23424 4483 24430
rect 4163 23360 4171 23424
rect 4235 23360 4251 23424
rect 4315 23360 4331 23424
rect 4395 23360 4411 23424
rect 4475 23360 4483 23424
rect 4163 22336 4483 23360
rect 4163 22272 4171 22336
rect 4235 22272 4251 22336
rect 4315 22272 4331 22336
rect 4395 22272 4411 22336
rect 4475 22272 4483 22336
rect 4163 21248 4483 22272
rect 4163 21184 4171 21248
rect 4235 21184 4251 21248
rect 4315 21184 4331 21248
rect 4395 21184 4411 21248
rect 4475 21184 4483 21248
rect 4163 20160 4483 21184
rect 4163 20096 4171 20160
rect 4235 20096 4251 20160
rect 4315 20096 4331 20160
rect 4395 20096 4411 20160
rect 4475 20096 4483 20160
rect 4163 19072 4483 20096
rect 4163 19008 4171 19072
rect 4235 19008 4251 19072
rect 4315 19008 4331 19072
rect 4395 19008 4411 19072
rect 4475 19008 4483 19072
rect 4163 18274 4483 19008
rect 4163 18038 4205 18274
rect 4441 18038 4483 18274
rect 4163 17984 4483 18038
rect 4163 17920 4171 17984
rect 4235 17920 4251 17984
rect 4315 17920 4331 17984
rect 4395 17920 4411 17984
rect 4475 17920 4483 17984
rect 4163 16896 4483 17920
rect 4163 16832 4171 16896
rect 4235 16832 4251 16896
rect 4315 16832 4331 16896
rect 4395 16832 4411 16896
rect 4475 16832 4483 16896
rect 4163 15808 4483 16832
rect 4163 15744 4171 15808
rect 4235 15744 4251 15808
rect 4315 15744 4331 15808
rect 4395 15744 4411 15808
rect 4475 15744 4483 15808
rect 4163 14720 4483 15744
rect 4163 14656 4171 14720
rect 4235 14656 4251 14720
rect 4315 14656 4331 14720
rect 4395 14656 4411 14720
rect 4475 14656 4483 14720
rect 4163 13632 4483 14656
rect 4163 13568 4171 13632
rect 4235 13568 4251 13632
rect 4315 13568 4331 13632
rect 4395 13568 4411 13632
rect 4475 13568 4483 13632
rect 4163 12544 4483 13568
rect 4163 12480 4171 12544
rect 4235 12480 4251 12544
rect 4315 12480 4331 12544
rect 4395 12480 4411 12544
rect 4475 12480 4483 12544
rect 4163 11882 4483 12480
rect 4163 11646 4205 11882
rect 4441 11646 4483 11882
rect 4163 11456 4483 11646
rect 4163 11392 4171 11456
rect 4235 11392 4251 11456
rect 4315 11392 4331 11456
rect 4395 11392 4411 11456
rect 4475 11392 4483 11456
rect 4163 10368 4483 11392
rect 4163 10304 4171 10368
rect 4235 10304 4251 10368
rect 4315 10304 4331 10368
rect 4395 10304 4411 10368
rect 4475 10304 4483 10368
rect 4163 9280 4483 10304
rect 4163 9216 4171 9280
rect 4235 9216 4251 9280
rect 4315 9216 4331 9280
rect 4395 9216 4411 9280
rect 4475 9216 4483 9280
rect 4163 8192 4483 9216
rect 4163 8128 4171 8192
rect 4235 8128 4251 8192
rect 4315 8128 4331 8192
rect 4395 8128 4411 8192
rect 4475 8128 4483 8192
rect 4163 7104 4483 8128
rect 4163 7040 4171 7104
rect 4235 7040 4251 7104
rect 4315 7040 4331 7104
rect 4395 7040 4411 7104
rect 4475 7040 4483 7104
rect 4163 6016 4483 7040
rect 4163 5952 4171 6016
rect 4235 5952 4251 6016
rect 4315 5952 4331 6016
rect 4395 5952 4411 6016
rect 4475 5952 4483 6016
rect 4163 5490 4483 5952
rect 4163 5254 4205 5490
rect 4441 5254 4483 5490
rect 4163 4928 4483 5254
rect 4163 4864 4171 4928
rect 4235 4864 4251 4928
rect 4315 4864 4331 4928
rect 4395 4864 4411 4928
rect 4475 4864 4483 4928
rect 4163 3840 4483 4864
rect 4163 3776 4171 3840
rect 4235 3776 4251 3840
rect 4315 3776 4331 3840
rect 4395 3776 4411 3840
rect 4475 3776 4483 3840
rect 4163 2752 4483 3776
rect 4163 2688 4171 2752
rect 4235 2688 4251 2752
rect 4315 2688 4331 2752
rect 4395 2688 4411 2752
rect 4475 2688 4483 2752
rect 4163 2128 4483 2688
rect 4823 27232 5143 27792
rect 4823 27168 4831 27232
rect 4895 27168 4911 27232
rect 4975 27168 4991 27232
rect 5055 27168 5071 27232
rect 5135 27168 5143 27232
rect 4823 26144 5143 27168
rect 4823 26080 4831 26144
rect 4895 26080 4911 26144
rect 4975 26080 4991 26144
rect 5055 26080 5071 26144
rect 5135 26080 5143 26144
rect 4823 25326 5143 26080
rect 4823 25090 4865 25326
rect 5101 25090 5143 25326
rect 4823 25056 5143 25090
rect 4823 24992 4831 25056
rect 4895 24992 4911 25056
rect 4975 24992 4991 25056
rect 5055 24992 5071 25056
rect 5135 24992 5143 25056
rect 4823 23968 5143 24992
rect 4823 23904 4831 23968
rect 4895 23904 4911 23968
rect 4975 23904 4991 23968
rect 5055 23904 5071 23968
rect 5135 23904 5143 23968
rect 4823 22880 5143 23904
rect 4823 22816 4831 22880
rect 4895 22816 4911 22880
rect 4975 22816 4991 22880
rect 5055 22816 5071 22880
rect 5135 22816 5143 22880
rect 4823 21792 5143 22816
rect 4823 21728 4831 21792
rect 4895 21728 4911 21792
rect 4975 21728 4991 21792
rect 5055 21728 5071 21792
rect 5135 21728 5143 21792
rect 4823 20704 5143 21728
rect 4823 20640 4831 20704
rect 4895 20640 4911 20704
rect 4975 20640 4991 20704
rect 5055 20640 5071 20704
rect 5135 20640 5143 20704
rect 4823 19616 5143 20640
rect 4823 19552 4831 19616
rect 4895 19552 4911 19616
rect 4975 19552 4991 19616
rect 5055 19552 5071 19616
rect 5135 19552 5143 19616
rect 4823 18934 5143 19552
rect 4823 18698 4865 18934
rect 5101 18698 5143 18934
rect 4823 18528 5143 18698
rect 4823 18464 4831 18528
rect 4895 18464 4911 18528
rect 4975 18464 4991 18528
rect 5055 18464 5071 18528
rect 5135 18464 5143 18528
rect 4823 17440 5143 18464
rect 4823 17376 4831 17440
rect 4895 17376 4911 17440
rect 4975 17376 4991 17440
rect 5055 17376 5071 17440
rect 5135 17376 5143 17440
rect 4823 16352 5143 17376
rect 4823 16288 4831 16352
rect 4895 16288 4911 16352
rect 4975 16288 4991 16352
rect 5055 16288 5071 16352
rect 5135 16288 5143 16352
rect 4823 15264 5143 16288
rect 4823 15200 4831 15264
rect 4895 15200 4911 15264
rect 4975 15200 4991 15264
rect 5055 15200 5071 15264
rect 5135 15200 5143 15264
rect 4823 14176 5143 15200
rect 4823 14112 4831 14176
rect 4895 14112 4911 14176
rect 4975 14112 4991 14176
rect 5055 14112 5071 14176
rect 5135 14112 5143 14176
rect 4823 13088 5143 14112
rect 4823 13024 4831 13088
rect 4895 13024 4911 13088
rect 4975 13024 4991 13088
rect 5055 13024 5071 13088
rect 5135 13024 5143 13088
rect 4823 12542 5143 13024
rect 4823 12306 4865 12542
rect 5101 12306 5143 12542
rect 4823 12000 5143 12306
rect 4823 11936 4831 12000
rect 4895 11936 4911 12000
rect 4975 11936 4991 12000
rect 5055 11936 5071 12000
rect 5135 11936 5143 12000
rect 4823 10912 5143 11936
rect 4823 10848 4831 10912
rect 4895 10848 4911 10912
rect 4975 10848 4991 10912
rect 5055 10848 5071 10912
rect 5135 10848 5143 10912
rect 4823 9824 5143 10848
rect 4823 9760 4831 9824
rect 4895 9760 4911 9824
rect 4975 9760 4991 9824
rect 5055 9760 5071 9824
rect 5135 9760 5143 9824
rect 4823 8736 5143 9760
rect 4823 8672 4831 8736
rect 4895 8672 4911 8736
rect 4975 8672 4991 8736
rect 5055 8672 5071 8736
rect 5135 8672 5143 8736
rect 4823 7648 5143 8672
rect 4823 7584 4831 7648
rect 4895 7584 4911 7648
rect 4975 7584 4991 7648
rect 5055 7584 5071 7648
rect 5135 7584 5143 7648
rect 4823 6560 5143 7584
rect 4823 6496 4831 6560
rect 4895 6496 4911 6560
rect 4975 6496 4991 6560
rect 5055 6496 5071 6560
rect 5135 6496 5143 6560
rect 4823 6150 5143 6496
rect 4823 5914 4865 6150
rect 5101 5914 5143 6150
rect 4823 5472 5143 5914
rect 4823 5408 4831 5472
rect 4895 5408 4911 5472
rect 4975 5408 4991 5472
rect 5055 5408 5071 5472
rect 5135 5408 5143 5472
rect 4823 4384 5143 5408
rect 4823 4320 4831 4384
rect 4895 4320 4911 4384
rect 4975 4320 4991 4384
rect 5055 4320 5071 4384
rect 5135 4320 5143 4384
rect 4823 3296 5143 4320
rect 4823 3232 4831 3296
rect 4895 3232 4911 3296
rect 4975 3232 4991 3296
rect 5055 3232 5071 3296
rect 5135 3232 5143 3296
rect 4823 2208 5143 3232
rect 4823 2144 4831 2208
rect 4895 2144 4911 2208
rect 4975 2144 4991 2208
rect 5055 2144 5071 2208
rect 5135 2144 5143 2208
rect 4823 2128 5143 2144
rect 10602 27776 10922 27792
rect 10602 27712 10610 27776
rect 10674 27712 10690 27776
rect 10754 27712 10770 27776
rect 10834 27712 10850 27776
rect 10914 27712 10922 27776
rect 10602 26688 10922 27712
rect 10602 26624 10610 26688
rect 10674 26624 10690 26688
rect 10754 26624 10770 26688
rect 10834 26624 10850 26688
rect 10914 26624 10922 26688
rect 10602 25600 10922 26624
rect 10602 25536 10610 25600
rect 10674 25536 10690 25600
rect 10754 25536 10770 25600
rect 10834 25536 10850 25600
rect 10914 25536 10922 25600
rect 10602 24666 10922 25536
rect 10602 24512 10644 24666
rect 10880 24512 10922 24666
rect 10602 24448 10610 24512
rect 10914 24448 10922 24512
rect 10602 24430 10644 24448
rect 10880 24430 10922 24448
rect 10602 23424 10922 24430
rect 10602 23360 10610 23424
rect 10674 23360 10690 23424
rect 10754 23360 10770 23424
rect 10834 23360 10850 23424
rect 10914 23360 10922 23424
rect 10602 22336 10922 23360
rect 10602 22272 10610 22336
rect 10674 22272 10690 22336
rect 10754 22272 10770 22336
rect 10834 22272 10850 22336
rect 10914 22272 10922 22336
rect 10602 21248 10922 22272
rect 10602 21184 10610 21248
rect 10674 21184 10690 21248
rect 10754 21184 10770 21248
rect 10834 21184 10850 21248
rect 10914 21184 10922 21248
rect 10602 20160 10922 21184
rect 10602 20096 10610 20160
rect 10674 20096 10690 20160
rect 10754 20096 10770 20160
rect 10834 20096 10850 20160
rect 10914 20096 10922 20160
rect 10602 19072 10922 20096
rect 10602 19008 10610 19072
rect 10674 19008 10690 19072
rect 10754 19008 10770 19072
rect 10834 19008 10850 19072
rect 10914 19008 10922 19072
rect 10602 18274 10922 19008
rect 10602 18038 10644 18274
rect 10880 18038 10922 18274
rect 10602 17984 10922 18038
rect 10602 17920 10610 17984
rect 10674 17920 10690 17984
rect 10754 17920 10770 17984
rect 10834 17920 10850 17984
rect 10914 17920 10922 17984
rect 10602 16896 10922 17920
rect 10602 16832 10610 16896
rect 10674 16832 10690 16896
rect 10754 16832 10770 16896
rect 10834 16832 10850 16896
rect 10914 16832 10922 16896
rect 10602 15808 10922 16832
rect 10602 15744 10610 15808
rect 10674 15744 10690 15808
rect 10754 15744 10770 15808
rect 10834 15744 10850 15808
rect 10914 15744 10922 15808
rect 10602 14720 10922 15744
rect 10602 14656 10610 14720
rect 10674 14656 10690 14720
rect 10754 14656 10770 14720
rect 10834 14656 10850 14720
rect 10914 14656 10922 14720
rect 10602 13632 10922 14656
rect 10602 13568 10610 13632
rect 10674 13568 10690 13632
rect 10754 13568 10770 13632
rect 10834 13568 10850 13632
rect 10914 13568 10922 13632
rect 10602 12544 10922 13568
rect 10602 12480 10610 12544
rect 10674 12480 10690 12544
rect 10754 12480 10770 12544
rect 10834 12480 10850 12544
rect 10914 12480 10922 12544
rect 10602 11882 10922 12480
rect 10602 11646 10644 11882
rect 10880 11646 10922 11882
rect 10602 11456 10922 11646
rect 10602 11392 10610 11456
rect 10674 11392 10690 11456
rect 10754 11392 10770 11456
rect 10834 11392 10850 11456
rect 10914 11392 10922 11456
rect 10602 10368 10922 11392
rect 10602 10304 10610 10368
rect 10674 10304 10690 10368
rect 10754 10304 10770 10368
rect 10834 10304 10850 10368
rect 10914 10304 10922 10368
rect 10602 9280 10922 10304
rect 10602 9216 10610 9280
rect 10674 9216 10690 9280
rect 10754 9216 10770 9280
rect 10834 9216 10850 9280
rect 10914 9216 10922 9280
rect 10602 8192 10922 9216
rect 10602 8128 10610 8192
rect 10674 8128 10690 8192
rect 10754 8128 10770 8192
rect 10834 8128 10850 8192
rect 10914 8128 10922 8192
rect 10602 7104 10922 8128
rect 10602 7040 10610 7104
rect 10674 7040 10690 7104
rect 10754 7040 10770 7104
rect 10834 7040 10850 7104
rect 10914 7040 10922 7104
rect 10602 6016 10922 7040
rect 10602 5952 10610 6016
rect 10674 5952 10690 6016
rect 10754 5952 10770 6016
rect 10834 5952 10850 6016
rect 10914 5952 10922 6016
rect 10602 5490 10922 5952
rect 10602 5254 10644 5490
rect 10880 5254 10922 5490
rect 10602 4928 10922 5254
rect 10602 4864 10610 4928
rect 10674 4864 10690 4928
rect 10754 4864 10770 4928
rect 10834 4864 10850 4928
rect 10914 4864 10922 4928
rect 10602 3840 10922 4864
rect 10602 3776 10610 3840
rect 10674 3776 10690 3840
rect 10754 3776 10770 3840
rect 10834 3776 10850 3840
rect 10914 3776 10922 3840
rect 10602 2752 10922 3776
rect 10602 2688 10610 2752
rect 10674 2688 10690 2752
rect 10754 2688 10770 2752
rect 10834 2688 10850 2752
rect 10914 2688 10922 2752
rect 10602 2128 10922 2688
rect 11262 27232 11582 27792
rect 11262 27168 11270 27232
rect 11334 27168 11350 27232
rect 11414 27168 11430 27232
rect 11494 27168 11510 27232
rect 11574 27168 11582 27232
rect 11262 26144 11582 27168
rect 11262 26080 11270 26144
rect 11334 26080 11350 26144
rect 11414 26080 11430 26144
rect 11494 26080 11510 26144
rect 11574 26080 11582 26144
rect 11262 25326 11582 26080
rect 11262 25090 11304 25326
rect 11540 25090 11582 25326
rect 11262 25056 11582 25090
rect 11262 24992 11270 25056
rect 11334 24992 11350 25056
rect 11414 24992 11430 25056
rect 11494 24992 11510 25056
rect 11574 24992 11582 25056
rect 11262 23968 11582 24992
rect 11262 23904 11270 23968
rect 11334 23904 11350 23968
rect 11414 23904 11430 23968
rect 11494 23904 11510 23968
rect 11574 23904 11582 23968
rect 11262 22880 11582 23904
rect 11262 22816 11270 22880
rect 11334 22816 11350 22880
rect 11414 22816 11430 22880
rect 11494 22816 11510 22880
rect 11574 22816 11582 22880
rect 11262 21792 11582 22816
rect 11262 21728 11270 21792
rect 11334 21728 11350 21792
rect 11414 21728 11430 21792
rect 11494 21728 11510 21792
rect 11574 21728 11582 21792
rect 11262 20704 11582 21728
rect 17041 27776 17361 27792
rect 17041 27712 17049 27776
rect 17113 27712 17129 27776
rect 17193 27712 17209 27776
rect 17273 27712 17289 27776
rect 17353 27712 17361 27776
rect 17041 26688 17361 27712
rect 17041 26624 17049 26688
rect 17113 26624 17129 26688
rect 17193 26624 17209 26688
rect 17273 26624 17289 26688
rect 17353 26624 17361 26688
rect 17041 25600 17361 26624
rect 17041 25536 17049 25600
rect 17113 25536 17129 25600
rect 17193 25536 17209 25600
rect 17273 25536 17289 25600
rect 17353 25536 17361 25600
rect 17041 24666 17361 25536
rect 17041 24512 17083 24666
rect 17319 24512 17361 24666
rect 17041 24448 17049 24512
rect 17353 24448 17361 24512
rect 17041 24430 17083 24448
rect 17319 24430 17361 24448
rect 17041 23424 17361 24430
rect 17041 23360 17049 23424
rect 17113 23360 17129 23424
rect 17193 23360 17209 23424
rect 17273 23360 17289 23424
rect 17353 23360 17361 23424
rect 17041 22336 17361 23360
rect 17041 22272 17049 22336
rect 17113 22272 17129 22336
rect 17193 22272 17209 22336
rect 17273 22272 17289 22336
rect 17353 22272 17361 22336
rect 17041 21248 17361 22272
rect 17041 21184 17049 21248
rect 17113 21184 17129 21248
rect 17193 21184 17209 21248
rect 17273 21184 17289 21248
rect 17353 21184 17361 21248
rect 15331 20772 15397 20773
rect 15331 20708 15332 20772
rect 15396 20708 15397 20772
rect 15331 20707 15397 20708
rect 11262 20640 11270 20704
rect 11334 20640 11350 20704
rect 11414 20640 11430 20704
rect 11494 20640 11510 20704
rect 11574 20640 11582 20704
rect 11262 19616 11582 20640
rect 11262 19552 11270 19616
rect 11334 19552 11350 19616
rect 11414 19552 11430 19616
rect 11494 19552 11510 19616
rect 11574 19552 11582 19616
rect 11262 18934 11582 19552
rect 11262 18698 11304 18934
rect 11540 18698 11582 18934
rect 11262 18528 11582 18698
rect 11262 18464 11270 18528
rect 11334 18464 11350 18528
rect 11414 18464 11430 18528
rect 11494 18464 11510 18528
rect 11574 18464 11582 18528
rect 11262 17440 11582 18464
rect 11262 17376 11270 17440
rect 11334 17376 11350 17440
rect 11414 17376 11430 17440
rect 11494 17376 11510 17440
rect 11574 17376 11582 17440
rect 11262 16352 11582 17376
rect 15334 17373 15394 20707
rect 15515 20500 15581 20501
rect 15515 20436 15516 20500
rect 15580 20436 15581 20500
rect 15515 20435 15581 20436
rect 15518 17917 15578 20435
rect 17041 20160 17361 21184
rect 17041 20096 17049 20160
rect 17113 20096 17129 20160
rect 17193 20096 17209 20160
rect 17273 20096 17289 20160
rect 17353 20096 17361 20160
rect 17041 19072 17361 20096
rect 17041 19008 17049 19072
rect 17113 19008 17129 19072
rect 17193 19008 17209 19072
rect 17273 19008 17289 19072
rect 17353 19008 17361 19072
rect 17041 18274 17361 19008
rect 17041 18038 17083 18274
rect 17319 18038 17361 18274
rect 17041 17984 17361 18038
rect 17041 17920 17049 17984
rect 17113 17920 17129 17984
rect 17193 17920 17209 17984
rect 17273 17920 17289 17984
rect 17353 17920 17361 17984
rect 15515 17916 15581 17917
rect 15515 17852 15516 17916
rect 15580 17852 15581 17916
rect 15515 17851 15581 17852
rect 15331 17372 15397 17373
rect 15331 17308 15332 17372
rect 15396 17308 15397 17372
rect 15331 17307 15397 17308
rect 11262 16288 11270 16352
rect 11334 16288 11350 16352
rect 11414 16288 11430 16352
rect 11494 16288 11510 16352
rect 11574 16288 11582 16352
rect 11262 15264 11582 16288
rect 11262 15200 11270 15264
rect 11334 15200 11350 15264
rect 11414 15200 11430 15264
rect 11494 15200 11510 15264
rect 11574 15200 11582 15264
rect 11262 14176 11582 15200
rect 11262 14112 11270 14176
rect 11334 14112 11350 14176
rect 11414 14112 11430 14176
rect 11494 14112 11510 14176
rect 11574 14112 11582 14176
rect 11262 13088 11582 14112
rect 11262 13024 11270 13088
rect 11334 13024 11350 13088
rect 11414 13024 11430 13088
rect 11494 13024 11510 13088
rect 11574 13024 11582 13088
rect 11262 12542 11582 13024
rect 11262 12306 11304 12542
rect 11540 12306 11582 12542
rect 11262 12000 11582 12306
rect 11262 11936 11270 12000
rect 11334 11936 11350 12000
rect 11414 11936 11430 12000
rect 11494 11936 11510 12000
rect 11574 11936 11582 12000
rect 11262 10912 11582 11936
rect 11262 10848 11270 10912
rect 11334 10848 11350 10912
rect 11414 10848 11430 10912
rect 11494 10848 11510 10912
rect 11574 10848 11582 10912
rect 11262 9824 11582 10848
rect 11262 9760 11270 9824
rect 11334 9760 11350 9824
rect 11414 9760 11430 9824
rect 11494 9760 11510 9824
rect 11574 9760 11582 9824
rect 11262 8736 11582 9760
rect 11262 8672 11270 8736
rect 11334 8672 11350 8736
rect 11414 8672 11430 8736
rect 11494 8672 11510 8736
rect 11574 8672 11582 8736
rect 11262 7648 11582 8672
rect 11262 7584 11270 7648
rect 11334 7584 11350 7648
rect 11414 7584 11430 7648
rect 11494 7584 11510 7648
rect 11574 7584 11582 7648
rect 11262 6560 11582 7584
rect 11262 6496 11270 6560
rect 11334 6496 11350 6560
rect 11414 6496 11430 6560
rect 11494 6496 11510 6560
rect 11574 6496 11582 6560
rect 11262 6150 11582 6496
rect 11262 5914 11304 6150
rect 11540 5914 11582 6150
rect 11262 5472 11582 5914
rect 11262 5408 11270 5472
rect 11334 5408 11350 5472
rect 11414 5408 11430 5472
rect 11494 5408 11510 5472
rect 11574 5408 11582 5472
rect 11262 4384 11582 5408
rect 11262 4320 11270 4384
rect 11334 4320 11350 4384
rect 11414 4320 11430 4384
rect 11494 4320 11510 4384
rect 11574 4320 11582 4384
rect 11262 3296 11582 4320
rect 11262 3232 11270 3296
rect 11334 3232 11350 3296
rect 11414 3232 11430 3296
rect 11494 3232 11510 3296
rect 11574 3232 11582 3296
rect 11262 2208 11582 3232
rect 11262 2144 11270 2208
rect 11334 2144 11350 2208
rect 11414 2144 11430 2208
rect 11494 2144 11510 2208
rect 11574 2144 11582 2208
rect 11262 2128 11582 2144
rect 17041 16896 17361 17920
rect 17041 16832 17049 16896
rect 17113 16832 17129 16896
rect 17193 16832 17209 16896
rect 17273 16832 17289 16896
rect 17353 16832 17361 16896
rect 17041 15808 17361 16832
rect 17041 15744 17049 15808
rect 17113 15744 17129 15808
rect 17193 15744 17209 15808
rect 17273 15744 17289 15808
rect 17353 15744 17361 15808
rect 17041 14720 17361 15744
rect 17041 14656 17049 14720
rect 17113 14656 17129 14720
rect 17193 14656 17209 14720
rect 17273 14656 17289 14720
rect 17353 14656 17361 14720
rect 17041 13632 17361 14656
rect 17041 13568 17049 13632
rect 17113 13568 17129 13632
rect 17193 13568 17209 13632
rect 17273 13568 17289 13632
rect 17353 13568 17361 13632
rect 17041 12544 17361 13568
rect 17041 12480 17049 12544
rect 17113 12480 17129 12544
rect 17193 12480 17209 12544
rect 17273 12480 17289 12544
rect 17353 12480 17361 12544
rect 17041 11882 17361 12480
rect 17041 11646 17083 11882
rect 17319 11646 17361 11882
rect 17041 11456 17361 11646
rect 17041 11392 17049 11456
rect 17113 11392 17129 11456
rect 17193 11392 17209 11456
rect 17273 11392 17289 11456
rect 17353 11392 17361 11456
rect 17041 10368 17361 11392
rect 17041 10304 17049 10368
rect 17113 10304 17129 10368
rect 17193 10304 17209 10368
rect 17273 10304 17289 10368
rect 17353 10304 17361 10368
rect 17041 9280 17361 10304
rect 17041 9216 17049 9280
rect 17113 9216 17129 9280
rect 17193 9216 17209 9280
rect 17273 9216 17289 9280
rect 17353 9216 17361 9280
rect 17041 8192 17361 9216
rect 17041 8128 17049 8192
rect 17113 8128 17129 8192
rect 17193 8128 17209 8192
rect 17273 8128 17289 8192
rect 17353 8128 17361 8192
rect 17041 7104 17361 8128
rect 17041 7040 17049 7104
rect 17113 7040 17129 7104
rect 17193 7040 17209 7104
rect 17273 7040 17289 7104
rect 17353 7040 17361 7104
rect 17041 6016 17361 7040
rect 17041 5952 17049 6016
rect 17113 5952 17129 6016
rect 17193 5952 17209 6016
rect 17273 5952 17289 6016
rect 17353 5952 17361 6016
rect 17041 5490 17361 5952
rect 17041 5254 17083 5490
rect 17319 5254 17361 5490
rect 17041 4928 17361 5254
rect 17041 4864 17049 4928
rect 17113 4864 17129 4928
rect 17193 4864 17209 4928
rect 17273 4864 17289 4928
rect 17353 4864 17361 4928
rect 17041 3840 17361 4864
rect 17041 3776 17049 3840
rect 17113 3776 17129 3840
rect 17193 3776 17209 3840
rect 17273 3776 17289 3840
rect 17353 3776 17361 3840
rect 17041 2752 17361 3776
rect 17041 2688 17049 2752
rect 17113 2688 17129 2752
rect 17193 2688 17209 2752
rect 17273 2688 17289 2752
rect 17353 2688 17361 2752
rect 17041 2128 17361 2688
rect 17701 27232 18021 27792
rect 17701 27168 17709 27232
rect 17773 27168 17789 27232
rect 17853 27168 17869 27232
rect 17933 27168 17949 27232
rect 18013 27168 18021 27232
rect 17701 26144 18021 27168
rect 17701 26080 17709 26144
rect 17773 26080 17789 26144
rect 17853 26080 17869 26144
rect 17933 26080 17949 26144
rect 18013 26080 18021 26144
rect 17701 25326 18021 26080
rect 17701 25090 17743 25326
rect 17979 25090 18021 25326
rect 17701 25056 18021 25090
rect 17701 24992 17709 25056
rect 17773 24992 17789 25056
rect 17853 24992 17869 25056
rect 17933 24992 17949 25056
rect 18013 24992 18021 25056
rect 17701 23968 18021 24992
rect 17701 23904 17709 23968
rect 17773 23904 17789 23968
rect 17853 23904 17869 23968
rect 17933 23904 17949 23968
rect 18013 23904 18021 23968
rect 17701 22880 18021 23904
rect 17701 22816 17709 22880
rect 17773 22816 17789 22880
rect 17853 22816 17869 22880
rect 17933 22816 17949 22880
rect 18013 22816 18021 22880
rect 17701 21792 18021 22816
rect 17701 21728 17709 21792
rect 17773 21728 17789 21792
rect 17853 21728 17869 21792
rect 17933 21728 17949 21792
rect 18013 21728 18021 21792
rect 17701 20704 18021 21728
rect 17701 20640 17709 20704
rect 17773 20640 17789 20704
rect 17853 20640 17869 20704
rect 17933 20640 17949 20704
rect 18013 20640 18021 20704
rect 17701 19616 18021 20640
rect 17701 19552 17709 19616
rect 17773 19552 17789 19616
rect 17853 19552 17869 19616
rect 17933 19552 17949 19616
rect 18013 19552 18021 19616
rect 17701 18934 18021 19552
rect 17701 18698 17743 18934
rect 17979 18698 18021 18934
rect 17701 18528 18021 18698
rect 17701 18464 17709 18528
rect 17773 18464 17789 18528
rect 17853 18464 17869 18528
rect 17933 18464 17949 18528
rect 18013 18464 18021 18528
rect 17701 17440 18021 18464
rect 17701 17376 17709 17440
rect 17773 17376 17789 17440
rect 17853 17376 17869 17440
rect 17933 17376 17949 17440
rect 18013 17376 18021 17440
rect 17701 16352 18021 17376
rect 17701 16288 17709 16352
rect 17773 16288 17789 16352
rect 17853 16288 17869 16352
rect 17933 16288 17949 16352
rect 18013 16288 18021 16352
rect 17701 15264 18021 16288
rect 17701 15200 17709 15264
rect 17773 15200 17789 15264
rect 17853 15200 17869 15264
rect 17933 15200 17949 15264
rect 18013 15200 18021 15264
rect 17701 14176 18021 15200
rect 17701 14112 17709 14176
rect 17773 14112 17789 14176
rect 17853 14112 17869 14176
rect 17933 14112 17949 14176
rect 18013 14112 18021 14176
rect 17701 13088 18021 14112
rect 17701 13024 17709 13088
rect 17773 13024 17789 13088
rect 17853 13024 17869 13088
rect 17933 13024 17949 13088
rect 18013 13024 18021 13088
rect 17701 12542 18021 13024
rect 17701 12306 17743 12542
rect 17979 12306 18021 12542
rect 17701 12000 18021 12306
rect 17701 11936 17709 12000
rect 17773 11936 17789 12000
rect 17853 11936 17869 12000
rect 17933 11936 17949 12000
rect 18013 11936 18021 12000
rect 17701 10912 18021 11936
rect 17701 10848 17709 10912
rect 17773 10848 17789 10912
rect 17853 10848 17869 10912
rect 17933 10848 17949 10912
rect 18013 10848 18021 10912
rect 17701 9824 18021 10848
rect 17701 9760 17709 9824
rect 17773 9760 17789 9824
rect 17853 9760 17869 9824
rect 17933 9760 17949 9824
rect 18013 9760 18021 9824
rect 17701 8736 18021 9760
rect 17701 8672 17709 8736
rect 17773 8672 17789 8736
rect 17853 8672 17869 8736
rect 17933 8672 17949 8736
rect 18013 8672 18021 8736
rect 17701 7648 18021 8672
rect 17701 7584 17709 7648
rect 17773 7584 17789 7648
rect 17853 7584 17869 7648
rect 17933 7584 17949 7648
rect 18013 7584 18021 7648
rect 17701 6560 18021 7584
rect 17701 6496 17709 6560
rect 17773 6496 17789 6560
rect 17853 6496 17869 6560
rect 17933 6496 17949 6560
rect 18013 6496 18021 6560
rect 17701 6150 18021 6496
rect 17701 5914 17743 6150
rect 17979 5914 18021 6150
rect 17701 5472 18021 5914
rect 17701 5408 17709 5472
rect 17773 5408 17789 5472
rect 17853 5408 17869 5472
rect 17933 5408 17949 5472
rect 18013 5408 18021 5472
rect 17701 4384 18021 5408
rect 17701 4320 17709 4384
rect 17773 4320 17789 4384
rect 17853 4320 17869 4384
rect 17933 4320 17949 4384
rect 18013 4320 18021 4384
rect 17701 3296 18021 4320
rect 17701 3232 17709 3296
rect 17773 3232 17789 3296
rect 17853 3232 17869 3296
rect 17933 3232 17949 3296
rect 18013 3232 18021 3296
rect 17701 2208 18021 3232
rect 17701 2144 17709 2208
rect 17773 2144 17789 2208
rect 17853 2144 17869 2208
rect 17933 2144 17949 2208
rect 18013 2144 18021 2208
rect 17701 2128 18021 2144
rect 23480 27776 23800 27792
rect 23480 27712 23488 27776
rect 23552 27712 23568 27776
rect 23632 27712 23648 27776
rect 23712 27712 23728 27776
rect 23792 27712 23800 27776
rect 23480 26688 23800 27712
rect 23480 26624 23488 26688
rect 23552 26624 23568 26688
rect 23632 26624 23648 26688
rect 23712 26624 23728 26688
rect 23792 26624 23800 26688
rect 23480 25600 23800 26624
rect 23480 25536 23488 25600
rect 23552 25536 23568 25600
rect 23632 25536 23648 25600
rect 23712 25536 23728 25600
rect 23792 25536 23800 25600
rect 23480 24666 23800 25536
rect 23480 24512 23522 24666
rect 23758 24512 23800 24666
rect 23480 24448 23488 24512
rect 23792 24448 23800 24512
rect 23480 24430 23522 24448
rect 23758 24430 23800 24448
rect 23480 23424 23800 24430
rect 23480 23360 23488 23424
rect 23552 23360 23568 23424
rect 23632 23360 23648 23424
rect 23712 23360 23728 23424
rect 23792 23360 23800 23424
rect 23480 22336 23800 23360
rect 23480 22272 23488 22336
rect 23552 22272 23568 22336
rect 23632 22272 23648 22336
rect 23712 22272 23728 22336
rect 23792 22272 23800 22336
rect 23480 21248 23800 22272
rect 23480 21184 23488 21248
rect 23552 21184 23568 21248
rect 23632 21184 23648 21248
rect 23712 21184 23728 21248
rect 23792 21184 23800 21248
rect 23480 20160 23800 21184
rect 23480 20096 23488 20160
rect 23552 20096 23568 20160
rect 23632 20096 23648 20160
rect 23712 20096 23728 20160
rect 23792 20096 23800 20160
rect 23480 19072 23800 20096
rect 23480 19008 23488 19072
rect 23552 19008 23568 19072
rect 23632 19008 23648 19072
rect 23712 19008 23728 19072
rect 23792 19008 23800 19072
rect 23480 18274 23800 19008
rect 23480 18038 23522 18274
rect 23758 18038 23800 18274
rect 23480 17984 23800 18038
rect 23480 17920 23488 17984
rect 23552 17920 23568 17984
rect 23632 17920 23648 17984
rect 23712 17920 23728 17984
rect 23792 17920 23800 17984
rect 23480 16896 23800 17920
rect 23480 16832 23488 16896
rect 23552 16832 23568 16896
rect 23632 16832 23648 16896
rect 23712 16832 23728 16896
rect 23792 16832 23800 16896
rect 23480 15808 23800 16832
rect 23480 15744 23488 15808
rect 23552 15744 23568 15808
rect 23632 15744 23648 15808
rect 23712 15744 23728 15808
rect 23792 15744 23800 15808
rect 23480 14720 23800 15744
rect 23480 14656 23488 14720
rect 23552 14656 23568 14720
rect 23632 14656 23648 14720
rect 23712 14656 23728 14720
rect 23792 14656 23800 14720
rect 23480 13632 23800 14656
rect 23480 13568 23488 13632
rect 23552 13568 23568 13632
rect 23632 13568 23648 13632
rect 23712 13568 23728 13632
rect 23792 13568 23800 13632
rect 23480 12544 23800 13568
rect 23480 12480 23488 12544
rect 23552 12480 23568 12544
rect 23632 12480 23648 12544
rect 23712 12480 23728 12544
rect 23792 12480 23800 12544
rect 23480 11882 23800 12480
rect 23480 11646 23522 11882
rect 23758 11646 23800 11882
rect 23480 11456 23800 11646
rect 23480 11392 23488 11456
rect 23552 11392 23568 11456
rect 23632 11392 23648 11456
rect 23712 11392 23728 11456
rect 23792 11392 23800 11456
rect 23480 10368 23800 11392
rect 23480 10304 23488 10368
rect 23552 10304 23568 10368
rect 23632 10304 23648 10368
rect 23712 10304 23728 10368
rect 23792 10304 23800 10368
rect 23480 9280 23800 10304
rect 23480 9216 23488 9280
rect 23552 9216 23568 9280
rect 23632 9216 23648 9280
rect 23712 9216 23728 9280
rect 23792 9216 23800 9280
rect 23480 8192 23800 9216
rect 23480 8128 23488 8192
rect 23552 8128 23568 8192
rect 23632 8128 23648 8192
rect 23712 8128 23728 8192
rect 23792 8128 23800 8192
rect 23480 7104 23800 8128
rect 23480 7040 23488 7104
rect 23552 7040 23568 7104
rect 23632 7040 23648 7104
rect 23712 7040 23728 7104
rect 23792 7040 23800 7104
rect 23480 6016 23800 7040
rect 23480 5952 23488 6016
rect 23552 5952 23568 6016
rect 23632 5952 23648 6016
rect 23712 5952 23728 6016
rect 23792 5952 23800 6016
rect 23480 5490 23800 5952
rect 23480 5254 23522 5490
rect 23758 5254 23800 5490
rect 23480 4928 23800 5254
rect 23480 4864 23488 4928
rect 23552 4864 23568 4928
rect 23632 4864 23648 4928
rect 23712 4864 23728 4928
rect 23792 4864 23800 4928
rect 23480 3840 23800 4864
rect 23480 3776 23488 3840
rect 23552 3776 23568 3840
rect 23632 3776 23648 3840
rect 23712 3776 23728 3840
rect 23792 3776 23800 3840
rect 23480 2752 23800 3776
rect 23480 2688 23488 2752
rect 23552 2688 23568 2752
rect 23632 2688 23648 2752
rect 23712 2688 23728 2752
rect 23792 2688 23800 2752
rect 23480 2128 23800 2688
rect 24140 27232 24460 27792
rect 24140 27168 24148 27232
rect 24212 27168 24228 27232
rect 24292 27168 24308 27232
rect 24372 27168 24388 27232
rect 24452 27168 24460 27232
rect 24140 26144 24460 27168
rect 24140 26080 24148 26144
rect 24212 26080 24228 26144
rect 24292 26080 24308 26144
rect 24372 26080 24388 26144
rect 24452 26080 24460 26144
rect 24140 25326 24460 26080
rect 24140 25090 24182 25326
rect 24418 25090 24460 25326
rect 24140 25056 24460 25090
rect 24140 24992 24148 25056
rect 24212 24992 24228 25056
rect 24292 24992 24308 25056
rect 24372 24992 24388 25056
rect 24452 24992 24460 25056
rect 24140 23968 24460 24992
rect 24140 23904 24148 23968
rect 24212 23904 24228 23968
rect 24292 23904 24308 23968
rect 24372 23904 24388 23968
rect 24452 23904 24460 23968
rect 24140 22880 24460 23904
rect 24140 22816 24148 22880
rect 24212 22816 24228 22880
rect 24292 22816 24308 22880
rect 24372 22816 24388 22880
rect 24452 22816 24460 22880
rect 24140 21792 24460 22816
rect 24140 21728 24148 21792
rect 24212 21728 24228 21792
rect 24292 21728 24308 21792
rect 24372 21728 24388 21792
rect 24452 21728 24460 21792
rect 24140 20704 24460 21728
rect 24140 20640 24148 20704
rect 24212 20640 24228 20704
rect 24292 20640 24308 20704
rect 24372 20640 24388 20704
rect 24452 20640 24460 20704
rect 24140 19616 24460 20640
rect 24140 19552 24148 19616
rect 24212 19552 24228 19616
rect 24292 19552 24308 19616
rect 24372 19552 24388 19616
rect 24452 19552 24460 19616
rect 24140 18934 24460 19552
rect 24140 18698 24182 18934
rect 24418 18698 24460 18934
rect 24140 18528 24460 18698
rect 24140 18464 24148 18528
rect 24212 18464 24228 18528
rect 24292 18464 24308 18528
rect 24372 18464 24388 18528
rect 24452 18464 24460 18528
rect 24140 17440 24460 18464
rect 24140 17376 24148 17440
rect 24212 17376 24228 17440
rect 24292 17376 24308 17440
rect 24372 17376 24388 17440
rect 24452 17376 24460 17440
rect 24140 16352 24460 17376
rect 24140 16288 24148 16352
rect 24212 16288 24228 16352
rect 24292 16288 24308 16352
rect 24372 16288 24388 16352
rect 24452 16288 24460 16352
rect 24140 15264 24460 16288
rect 24140 15200 24148 15264
rect 24212 15200 24228 15264
rect 24292 15200 24308 15264
rect 24372 15200 24388 15264
rect 24452 15200 24460 15264
rect 24140 14176 24460 15200
rect 24140 14112 24148 14176
rect 24212 14112 24228 14176
rect 24292 14112 24308 14176
rect 24372 14112 24388 14176
rect 24452 14112 24460 14176
rect 24140 13088 24460 14112
rect 24140 13024 24148 13088
rect 24212 13024 24228 13088
rect 24292 13024 24308 13088
rect 24372 13024 24388 13088
rect 24452 13024 24460 13088
rect 24140 12542 24460 13024
rect 24140 12306 24182 12542
rect 24418 12306 24460 12542
rect 24140 12000 24460 12306
rect 24140 11936 24148 12000
rect 24212 11936 24228 12000
rect 24292 11936 24308 12000
rect 24372 11936 24388 12000
rect 24452 11936 24460 12000
rect 24140 10912 24460 11936
rect 24140 10848 24148 10912
rect 24212 10848 24228 10912
rect 24292 10848 24308 10912
rect 24372 10848 24388 10912
rect 24452 10848 24460 10912
rect 24140 9824 24460 10848
rect 24140 9760 24148 9824
rect 24212 9760 24228 9824
rect 24292 9760 24308 9824
rect 24372 9760 24388 9824
rect 24452 9760 24460 9824
rect 24140 8736 24460 9760
rect 24140 8672 24148 8736
rect 24212 8672 24228 8736
rect 24292 8672 24308 8736
rect 24372 8672 24388 8736
rect 24452 8672 24460 8736
rect 24140 7648 24460 8672
rect 24140 7584 24148 7648
rect 24212 7584 24228 7648
rect 24292 7584 24308 7648
rect 24372 7584 24388 7648
rect 24452 7584 24460 7648
rect 24140 6560 24460 7584
rect 24140 6496 24148 6560
rect 24212 6496 24228 6560
rect 24292 6496 24308 6560
rect 24372 6496 24388 6560
rect 24452 6496 24460 6560
rect 24140 6150 24460 6496
rect 24140 5914 24182 6150
rect 24418 5914 24460 6150
rect 24140 5472 24460 5914
rect 24140 5408 24148 5472
rect 24212 5408 24228 5472
rect 24292 5408 24308 5472
rect 24372 5408 24388 5472
rect 24452 5408 24460 5472
rect 24140 4384 24460 5408
rect 24140 4320 24148 4384
rect 24212 4320 24228 4384
rect 24292 4320 24308 4384
rect 24372 4320 24388 4384
rect 24452 4320 24460 4384
rect 24140 3296 24460 4320
rect 24140 3232 24148 3296
rect 24212 3232 24228 3296
rect 24292 3232 24308 3296
rect 24372 3232 24388 3296
rect 24452 3232 24460 3296
rect 24140 2208 24460 3232
rect 24140 2144 24148 2208
rect 24212 2144 24228 2208
rect 24292 2144 24308 2208
rect 24372 2144 24388 2208
rect 24452 2144 24460 2208
rect 24140 2128 24460 2144
<< via4 >>
rect 4205 24512 4441 24666
rect 4205 24448 4235 24512
rect 4235 24448 4251 24512
rect 4251 24448 4315 24512
rect 4315 24448 4331 24512
rect 4331 24448 4395 24512
rect 4395 24448 4411 24512
rect 4411 24448 4441 24512
rect 4205 24430 4441 24448
rect 4205 18038 4441 18274
rect 4205 11646 4441 11882
rect 4205 5254 4441 5490
rect 4865 25090 5101 25326
rect 4865 18698 5101 18934
rect 4865 12306 5101 12542
rect 4865 5914 5101 6150
rect 10644 24512 10880 24666
rect 10644 24448 10674 24512
rect 10674 24448 10690 24512
rect 10690 24448 10754 24512
rect 10754 24448 10770 24512
rect 10770 24448 10834 24512
rect 10834 24448 10850 24512
rect 10850 24448 10880 24512
rect 10644 24430 10880 24448
rect 10644 18038 10880 18274
rect 10644 11646 10880 11882
rect 10644 5254 10880 5490
rect 11304 25090 11540 25326
rect 17083 24512 17319 24666
rect 17083 24448 17113 24512
rect 17113 24448 17129 24512
rect 17129 24448 17193 24512
rect 17193 24448 17209 24512
rect 17209 24448 17273 24512
rect 17273 24448 17289 24512
rect 17289 24448 17319 24512
rect 17083 24430 17319 24448
rect 11304 18698 11540 18934
rect 17083 18038 17319 18274
rect 11304 12306 11540 12542
rect 11304 5914 11540 6150
rect 17083 11646 17319 11882
rect 17083 5254 17319 5490
rect 17743 25090 17979 25326
rect 17743 18698 17979 18934
rect 17743 12306 17979 12542
rect 17743 5914 17979 6150
rect 23522 24512 23758 24666
rect 23522 24448 23552 24512
rect 23552 24448 23568 24512
rect 23568 24448 23632 24512
rect 23632 24448 23648 24512
rect 23648 24448 23712 24512
rect 23712 24448 23728 24512
rect 23728 24448 23758 24512
rect 23522 24430 23758 24448
rect 23522 18038 23758 18274
rect 23522 11646 23758 11882
rect 23522 5254 23758 5490
rect 24182 25090 24418 25326
rect 24182 18698 24418 18934
rect 24182 12306 24418 12542
rect 24182 5914 24418 6150
<< metal5 >>
rect 1056 25326 26912 25368
rect 1056 25090 4865 25326
rect 5101 25090 11304 25326
rect 11540 25090 17743 25326
rect 17979 25090 24182 25326
rect 24418 25090 26912 25326
rect 1056 25048 26912 25090
rect 1056 24666 26912 24708
rect 1056 24430 4205 24666
rect 4441 24430 10644 24666
rect 10880 24430 17083 24666
rect 17319 24430 23522 24666
rect 23758 24430 26912 24666
rect 1056 24388 26912 24430
rect 1056 18934 26912 18976
rect 1056 18698 4865 18934
rect 5101 18698 11304 18934
rect 11540 18698 17743 18934
rect 17979 18698 24182 18934
rect 24418 18698 26912 18934
rect 1056 18656 26912 18698
rect 1056 18274 26912 18316
rect 1056 18038 4205 18274
rect 4441 18038 10644 18274
rect 10880 18038 17083 18274
rect 17319 18038 23522 18274
rect 23758 18038 26912 18274
rect 1056 17996 26912 18038
rect 1056 12542 26912 12584
rect 1056 12306 4865 12542
rect 5101 12306 11304 12542
rect 11540 12306 17743 12542
rect 17979 12306 24182 12542
rect 24418 12306 26912 12542
rect 1056 12264 26912 12306
rect 1056 11882 26912 11924
rect 1056 11646 4205 11882
rect 4441 11646 10644 11882
rect 10880 11646 17083 11882
rect 17319 11646 23522 11882
rect 23758 11646 26912 11882
rect 1056 11604 26912 11646
rect 1056 6150 26912 6192
rect 1056 5914 4865 6150
rect 5101 5914 11304 6150
rect 11540 5914 17743 6150
rect 17979 5914 24182 6150
rect 24418 5914 26912 6150
rect 1056 5872 26912 5914
rect 1056 5490 26912 5532
rect 1056 5254 4205 5490
rect 4441 5254 10644 5490
rect 10880 5254 17083 5490
rect 17319 5254 23522 5490
rect 23758 5254 26912 5490
rect 1056 5212 26912 5254
use sky130_fd_sc_hd__buf_2  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17940 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14812 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15640 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0639_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0640_
timestamp 1698431365
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17480 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16468 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0646_
timestamp 1698431365
transform -1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0647_
timestamp 1698431365
transform -1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0648_
timestamp 1698431365
transform 1 0 17480 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17572 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1698431365
transform -1 0 18768 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 19136 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1698431365
transform 1 0 17204 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0653_
timestamp 1698431365
transform -1 0 18676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 1698431365
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 18492 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0657_
timestamp 1698431365
transform -1 0 18400 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1698431365
transform -1 0 18492 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1698431365
transform -1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19596 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0661_
timestamp 1698431365
transform 1 0 18400 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0662_
timestamp 1698431365
transform 1 0 18492 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1698431365
transform -1 0 18768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 18768 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0665_
timestamp 1698431365
transform 1 0 17572 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1698431365
transform -1 0 17572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0667_
timestamp 1698431365
transform -1 0 18400 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0668_
timestamp 1698431365
transform -1 0 16744 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1698431365
transform -1 0 16376 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1698431365
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1698431365
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0672_
timestamp 1698431365
transform -1 0 17480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1698431365
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1698431365
transform -1 0 13156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0675_
timestamp 1698431365
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0676_
timestamp 1698431365
transform -1 0 16008 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1698431365
transform -1 0 15180 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1698431365
transform -1 0 15732 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0679_
timestamp 1698431365
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1698431365
transform 1 0 14168 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1698431365
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0682_
timestamp 1698431365
transform 1 0 13432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0683_
timestamp 1698431365
transform -1 0 17388 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1698431365
transform 1 0 13616 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1698431365
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0686_
timestamp 1698431365
transform -1 0 18676 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1698431365
transform 1 0 17940 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1698431365
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0689_
timestamp 1698431365
transform 1 0 19228 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1698431365
transform -1 0 20056 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1698431365
transform 1 0 20056 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0692_
timestamp 1698431365
transform 1 0 18124 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1698431365
transform 1 0 18952 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1698431365
transform -1 0 19136 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1698431365
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1698431365
transform -1 0 17940 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1698431365
transform -1 0 17940 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0698_
timestamp 1698431365
transform -1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0699_
timestamp 1698431365
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0700_
timestamp 1698431365
transform -1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1698431365
transform 1 0 11868 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1698431365
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0703_
timestamp 1698431365
transform -1 0 16008 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1698431365
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0705_
timestamp 1698431365
transform -1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17112 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1698431365
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0708_
timestamp 1698431365
transform 1 0 12604 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0709_
timestamp 1698431365
transform -1 0 15180 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1698431365
transform 1 0 12328 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1698431365
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1698431365
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0713_
timestamp 1698431365
transform -1 0 15640 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1698431365
transform 1 0 13708 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0715_
timestamp 1698431365
transform 1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 19044 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1698431365
transform -1 0 20148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19228 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1698431365
transform -1 0 20976 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0720_
timestamp 1698431365
transform -1 0 20332 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0721_
timestamp 1698431365
transform 1 0 19228 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 21620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1698431365
transform -1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0724_
timestamp 1698431365
transform 1 0 20608 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1698431365
transform 1 0 20516 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 21712 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0727_
timestamp 1698431365
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0728_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 21896 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0729_
timestamp 1698431365
transform 1 0 20884 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1698431365
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 20976 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1698431365
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1698431365
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0737_
timestamp 1698431365
transform 1 0 19228 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0738_
timestamp 1698431365
transform -1 0 20148 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0739_
timestamp 1698431365
transform 1 0 20148 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 1698431365
transform 1 0 18308 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0741_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0742_
timestamp 1698431365
transform -1 0 18768 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0743_
timestamp 1698431365
transform -1 0 19872 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0744_
timestamp 1698431365
transform -1 0 13984 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1698431365
transform 1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0746_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12144 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1698431365
transform -1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1698431365
transform -1 0 13984 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1698431365
transform -1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0750_
timestamp 1698431365
transform -1 0 13984 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0751_
timestamp 1698431365
transform 1 0 12972 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0752_
timestamp 1698431365
transform -1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 1698431365
transform -1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0754_
timestamp 1698431365
transform 1 0 15088 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0755_
timestamp 1698431365
transform -1 0 15916 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0756_
timestamp 1698431365
transform -1 0 16376 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0757_
timestamp 1698431365
transform 1 0 15548 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0758_
timestamp 1698431365
transform 1 0 14996 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1698431365
transform 1 0 15732 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0760_
timestamp 1698431365
transform 1 0 16192 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0761_
timestamp 1698431365
transform -1 0 14628 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0762_
timestamp 1698431365
transform -1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1698431365
transform -1 0 13248 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0764_
timestamp 1698431365
transform 1 0 14076 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0765_
timestamp 1698431365
transform -1 0 13524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1698431365
transform -1 0 13984 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0767_
timestamp 1698431365
transform -1 0 12972 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1698431365
transform -1 0 12328 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 1698431365
transform 1 0 10856 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0770_
timestamp 1698431365
transform 1 0 11592 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0771_
timestamp 1698431365
transform 1 0 11500 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1698431365
transform -1 0 11408 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0773_
timestamp 1698431365
transform -1 0 7728 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1698431365
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0775_
timestamp 1698431365
transform 1 0 4416 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0776_
timestamp 1698431365
transform -1 0 7728 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0777_
timestamp 1698431365
transform -1 0 7360 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0778_
timestamp 1698431365
transform -1 0 4876 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 1698431365
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1698431365
transform 1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 1698431365
transform 1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0782_
timestamp 1698431365
transform -1 0 7176 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0783_
timestamp 1698431365
transform -1 0 4508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0784_
timestamp 1698431365
transform -1 0 3680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0785_
timestamp 1698431365
transform -1 0 7268 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0786_
timestamp 1698431365
transform 1 0 6256 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0787_
timestamp 1698431365
transform 1 0 7176 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0788_
timestamp 1698431365
transform 1 0 6532 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0789_
timestamp 1698431365
transform 1 0 6808 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1698431365
transform -1 0 6256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1698431365
transform -1 0 6900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0792_
timestamp 1698431365
transform 1 0 7728 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1698431365
transform 1 0 6256 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1698431365
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1698431365
transform 1 0 4968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0796_
timestamp 1698431365
transform -1 0 4968 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0797_
timestamp 1698431365
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0798_
timestamp 1698431365
transform 1 0 3772 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3680 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0800_
timestamp 1698431365
transform -1 0 4508 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0801_
timestamp 1698431365
transform 1 0 5152 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0802_
timestamp 1698431365
transform -1 0 6992 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1698431365
transform 1 0 5152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0804_
timestamp 1698431365
transform 1 0 3864 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0805_
timestamp 1698431365
transform -1 0 5612 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0806_
timestamp 1698431365
transform -1 0 5428 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0807_
timestamp 1698431365
transform -1 0 4876 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0808_
timestamp 1698431365
transform -1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1698431365
transform -1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0810_
timestamp 1698431365
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 1698431365
transform -1 0 5060 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0812_
timestamp 1698431365
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0813_
timestamp 1698431365
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 1698431365
transform 1 0 4416 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0815_
timestamp 1698431365
transform 1 0 4508 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0816_
timestamp 1698431365
transform 1 0 5704 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0817_
timestamp 1698431365
transform 1 0 5060 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0818_
timestamp 1698431365
transform -1 0 5980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 1698431365
transform 1 0 5520 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1698431365
transform 1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0821_
timestamp 1698431365
transform 1 0 5612 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0822_
timestamp 1698431365
transform -1 0 5244 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0823_
timestamp 1698431365
transform 1 0 4968 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0824_
timestamp 1698431365
transform -1 0 4876 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0825_
timestamp 1698431365
transform 1 0 3680 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0826_
timestamp 1698431365
transform 1 0 2852 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0827_
timestamp 1698431365
transform -1 0 4232 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0828_
timestamp 1698431365
transform 1 0 3772 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0829_
timestamp 1698431365
transform 1 0 2944 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0830_
timestamp 1698431365
transform -1 0 7636 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1698431365
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0832_
timestamp 1698431365
transform 1 0 5428 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0833_
timestamp 1698431365
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0834_
timestamp 1698431365
transform -1 0 6256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1698431365
transform -1 0 5428 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0836_
timestamp 1698431365
transform -1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1698431365
transform -1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1698431365
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0839_
timestamp 1698431365
transform -1 0 5796 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0840_
timestamp 1698431365
transform -1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1698431365
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0842_
timestamp 1698431365
transform -1 0 7636 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0843_
timestamp 1698431365
transform -1 0 6256 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0844_
timestamp 1698431365
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0845_
timestamp 1698431365
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0846_
timestamp 1698431365
transform -1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0847_
timestamp 1698431365
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1698431365
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0849_
timestamp 1698431365
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1698431365
transform -1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0851_
timestamp 1698431365
transform 1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0852_
timestamp 1698431365
transform -1 0 5428 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1698431365
transform -1 0 5704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0854_
timestamp 1698431365
transform -1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0855_
timestamp 1698431365
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0856_
timestamp 1698431365
transform 1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0857_
timestamp 1698431365
transform 1 0 3864 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0858_
timestamp 1698431365
transform 1 0 13800 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1698431365
transform -1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0860_
timestamp 1698431365
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0861_
timestamp 1698431365
transform -1 0 13248 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0862_
timestamp 1698431365
transform 1 0 13524 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0863_
timestamp 1698431365
transform -1 0 15272 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0864_
timestamp 1698431365
transform -1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1698431365
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0866_
timestamp 1698431365
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0867_
timestamp 1698431365
transform -1 0 12604 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1698431365
transform -1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1698431365
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0870_
timestamp 1698431365
transform 1 0 12512 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0871_
timestamp 1698431365
transform 1 0 12604 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1698431365
transform 1 0 13248 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1698431365
transform 1 0 13156 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0874_
timestamp 1698431365
transform 1 0 13248 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1698431365
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1698431365
transform -1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1698431365
transform -1 0 15088 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0878_
timestamp 1698431365
transform 1 0 14720 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0879_
timestamp 1698431365
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0880_
timestamp 1698431365
transform 1 0 15272 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1698431365
transform 1 0 18032 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0882_
timestamp 1698431365
transform 1 0 16008 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0883_
timestamp 1698431365
transform -1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0884_
timestamp 1698431365
transform 1 0 18124 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0885_
timestamp 1698431365
transform 1 0 16652 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0886_
timestamp 1698431365
transform 1 0 16744 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1698431365
transform -1 0 19320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0888_
timestamp 1698431365
transform 1 0 18400 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0889_
timestamp 1698431365
transform 1 0 18676 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1698431365
transform -1 0 21712 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1698431365
transform 1 0 18676 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0892_
timestamp 1698431365
transform 1 0 19688 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1698431365
transform -1 0 16468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1698431365
transform -1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1698431365
transform -1 0 19964 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0896_
timestamp 1698431365
transform 1 0 19320 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0897_
timestamp 1698431365
transform 1 0 19136 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0898_
timestamp 1698431365
transform -1 0 21528 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0899_
timestamp 1698431365
transform 1 0 19964 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1698431365
transform 1 0 20516 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0901_
timestamp 1698431365
transform 1 0 20056 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0902_
timestamp 1698431365
transform 1 0 17388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0903_
timestamp 1698431365
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1698431365
transform -1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0905_
timestamp 1698431365
transform -1 0 20516 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1698431365
transform -1 0 21252 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0907_
timestamp 1698431365
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0908_
timestamp 1698431365
transform -1 0 18768 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1698431365
transform -1 0 18676 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0910_
timestamp 1698431365
transform 1 0 16836 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0911_
timestamp 1698431365
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0912_
timestamp 1698431365
transform 1 0 17756 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0913_
timestamp 1698431365
transform 1 0 17112 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0914_
timestamp 1698431365
transform -1 0 8464 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1698431365
transform 1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0916_
timestamp 1698431365
transform 1 0 4692 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1698431365
transform -1 0 7912 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0918_
timestamp 1698431365
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0919_
timestamp 1698431365
transform -1 0 6256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1698431365
transform -1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1698431365
transform -1 0 10212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1698431365
transform 1 0 8464 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1698431365
transform -1 0 6532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 1698431365
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0925_
timestamp 1698431365
transform 1 0 5336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0926_
timestamp 1698431365
transform 1 0 7084 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0927_
timestamp 1698431365
transform 1 0 6808 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1698431365
transform 1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0929_
timestamp 1698431365
transform 1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0930_
timestamp 1698431365
transform -1 0 9476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0931_
timestamp 1698431365
transform -1 0 8648 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1698431365
transform -1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0933_
timestamp 1698431365
transform 1 0 8280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1698431365
transform -1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0935_
timestamp 1698431365
transform 1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0936_
timestamp 1698431365
transform -1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1698431365
transform -1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0938_
timestamp 1698431365
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0939_
timestamp 1698431365
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0940_
timestamp 1698431365
transform -1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0941_
timestamp 1698431365
transform 1 0 4232 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _0943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3312 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1698431365
transform 1 0 12512 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1698431365
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12420 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14076 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0948_
timestamp 1698431365
transform -1 0 13524 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1698431365
transform -1 0 13524 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14168 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0952_
timestamp 1698431365
transform 1 0 12328 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1698431365
transform -1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0954_
timestamp 1698431365
transform 1 0 14720 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0955_
timestamp 1698431365
transform -1 0 14720 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1698431365
transform -1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0957_
timestamp 1698431365
transform -1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0958_
timestamp 1698431365
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1698431365
transform -1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 1698431365
transform -1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1698431365
transform 1 0 11224 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0962_
timestamp 1698431365
transform -1 0 11224 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _0963_
timestamp 1698431365
transform 1 0 13524 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1698431365
transform 1 0 13524 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1698431365
transform 1 0 15272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0966_
timestamp 1698431365
transform 1 0 13156 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0967_
timestamp 1698431365
transform 1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1698431365
transform 1 0 9568 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1698431365
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0970_
timestamp 1698431365
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1698431365
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1698431365
transform 1 0 17480 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1698431365
transform 1 0 16376 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1698431365
transform -1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1698431365
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0976_
timestamp 1698431365
transform 1 0 14444 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1698431365
transform 1 0 16652 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0980_
timestamp 1698431365
transform -1 0 16376 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1698431365
transform 1 0 15364 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1698431365
transform -1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15640 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15732 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_4  _0985_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17940 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1698431365
transform 1 0 15640 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1698431365
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_4  _0988_
timestamp 1698431365
transform -1 0 16560 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_4  _0989_
timestamp 1698431365
transform 1 0 15180 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_4  _0990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 2116 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 3312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0992_
timestamp 1698431365
transform 1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1698431365
transform -1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1698431365
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1698431365
transform 1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1698431365
transform -1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1698431365
transform -1 0 11408 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1698431365
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1698431365
transform 1 0 19872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1698431365
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1698431365
transform -1 0 19044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1698431365
transform 1 0 13064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1003_
timestamp 1698431365
transform 1 0 14996 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1698431365
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1698431365
transform -1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1698431365
transform -1 0 13984 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1698431365
transform -1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1698431365
transform -1 0 18952 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1698431365
transform 1 0 19964 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1698431365
transform 1 0 19504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1698431365
transform 1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1698431365
transform 1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1698431365
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1014_
timestamp 1698431365
transform 1 0 15824 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1698431365
transform -1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1698431365
transform -1 0 20516 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1698431365
transform -1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1698431365
transform -1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1698431365
transform -1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1698431365
transform -1 0 22632 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1021_
timestamp 1698431365
transform 1 0 22356 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1022_
timestamp 1698431365
transform -1 0 23184 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 22632 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1024_
timestamp 1698431365
transform 1 0 23184 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1025_
timestamp 1698431365
transform -1 0 24748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1026_
timestamp 1698431365
transform -1 0 25300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1027_
timestamp 1698431365
transform 1 0 23460 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1698431365
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 1698431365
transform 1 0 14260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1030_
timestamp 1698431365
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1698431365
transform 1 0 13248 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1032_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1033_
timestamp 1698431365
transform -1 0 9384 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp 1698431365
transform 1 0 7452 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1035_
timestamp 1698431365
transform -1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1698431365
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1037_
timestamp 1698431365
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1038_
timestamp 1698431365
transform -1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1039_
timestamp 1698431365
transform -1 0 9016 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1040_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 8740 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1041_
timestamp 1698431365
transform 1 0 7544 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1698431365
transform 1 0 8280 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1043_
timestamp 1698431365
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1698431365
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1045_
timestamp 1698431365
transform -1 0 13984 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1046_
timestamp 1698431365
transform -1 0 14076 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1047_
timestamp 1698431365
transform -1 0 13248 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 1698431365
transform 1 0 8556 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1050_
timestamp 1698431365
transform 1 0 10120 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1698431365
transform 1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1052_
timestamp 1698431365
transform -1 0 14260 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1053_
timestamp 1698431365
transform 1 0 12972 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1054_
timestamp 1698431365
transform -1 0 12788 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1698431365
transform -1 0 13892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1698431365
transform 1 0 7636 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1698431365
transform 1 0 9108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1058_
timestamp 1698431365
transform -1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1059_
timestamp 1698431365
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1060_
timestamp 1698431365
transform 1 0 9568 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1698431365
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9476 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1698431365
transform 1 0 8096 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1064_
timestamp 1698431365
transform -1 0 12604 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1065_
timestamp 1698431365
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1066_
timestamp 1698431365
transform 1 0 10764 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1698431365
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1698431365
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1069_
timestamp 1698431365
transform 1 0 11592 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 1698431365
transform 1 0 11500 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1071_
timestamp 1698431365
transform -1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1072_
timestamp 1698431365
transform -1 0 12604 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1073_
timestamp 1698431365
transform 1 0 10948 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1074_
timestamp 1698431365
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 1698431365
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1076_
timestamp 1698431365
transform 1 0 10304 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1077_
timestamp 1698431365
transform -1 0 9476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1078_
timestamp 1698431365
transform -1 0 10304 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1079_
timestamp 1698431365
transform -1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1080_
timestamp 1698431365
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1698431365
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1698431365
transform 1 0 22172 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1698431365
transform 1 0 17112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1698431365
transform 1 0 22632 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1698431365
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1698431365
transform -1 0 20148 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1698431365
transform 1 0 19504 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1698431365
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1698431365
transform -1 0 18124 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1090_
timestamp 1698431365
transform -1 0 6348 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1698431365
transform 1 0 14352 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1698431365
transform 1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1698431365
transform -1 0 16468 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1698431365
transform -1 0 14904 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1698431365
transform 1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1698431365
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1698431365
transform -1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1698431365
transform -1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1698431365
transform 1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1698431365
transform -1 0 9200 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1101_
timestamp 1698431365
transform 1 0 2760 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1698431365
transform 1 0 6992 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1698431365
transform -1 0 2944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1698431365
transform -1 0 3588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1698431365
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1698431365
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1698431365
transform -1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1698431365
transform 1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1698431365
transform -1 0 7268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1698431365
transform -1 0 2944 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1698431365
transform 1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1112_
timestamp 1698431365
transform -1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1698431365
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1698431365
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1698431365
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1698431365
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1698431365
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1698431365
transform -1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1698431365
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1698431365
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1698431365
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1698431365
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1123_
timestamp 1698431365
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1698431365
transform -1 0 14996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1698431365
transform -1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1698431365
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1698431365
transform -1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1698431365
transform 1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1698431365
transform -1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1698431365
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1698431365
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1698431365
transform -1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1698431365
transform 1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1698431365
transform 1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1698431365
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1698431365
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1698431365
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1698431365
transform -1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1698431365
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1698431365
transform -1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1698431365
transform -1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1142_
timestamp 1698431365
transform -1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1698431365
transform -1 0 12604 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1144_
timestamp 1698431365
transform -1 0 10396 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1145_
timestamp 1698431365
transform -1 0 12144 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1146_
timestamp 1698431365
transform 1 0 11224 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1147_
timestamp 1698431365
transform 1 0 10856 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 1698431365
transform 1 0 11500 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1149_
timestamp 1698431365
transform -1 0 12236 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1150_
timestamp 1698431365
transform -1 0 11408 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1151_
timestamp 1698431365
transform -1 0 11776 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1152_
timestamp 1698431365
transform 1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1698431365
transform -1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1154_
timestamp 1698431365
transform 1 0 8188 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1155_
timestamp 1698431365
transform -1 0 9660 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1156_
timestamp 1698431365
transform 1 0 12328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1157_
timestamp 1698431365
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9568 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1159_
timestamp 1698431365
transform 1 0 9752 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1160_
timestamp 1698431365
transform 1 0 13340 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1161_
timestamp 1698431365
transform -1 0 9476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1163_
timestamp 1698431365
transform 1 0 10672 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1164_
timestamp 1698431365
transform 1 0 10304 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1165_
timestamp 1698431365
transform 1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1166_
timestamp 1698431365
transform -1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1167_
timestamp 1698431365
transform 1 0 8372 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 1698431365
transform 1 0 8924 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1169_
timestamp 1698431365
transform -1 0 13340 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1170_
timestamp 1698431365
transform 1 0 9660 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1171_
timestamp 1698431365
transform -1 0 12328 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1172_
timestamp 1698431365
transform -1 0 10488 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1173_
timestamp 1698431365
transform -1 0 10856 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _1174_
timestamp 1698431365
transform -1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1175_
timestamp 1698431365
transform 1 0 10488 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1698431365
transform -1 0 10212 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1177_
timestamp 1698431365
transform -1 0 9752 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1178_
timestamp 1698431365
transform -1 0 9292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1179_
timestamp 1698431365
transform -1 0 10488 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1180_
timestamp 1698431365
transform -1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 1698431365
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _1182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9752 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1183_
timestamp 1698431365
transform 1 0 9016 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_4  _1184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 10304 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1698431365
transform 1 0 7636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1698431365
transform 1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1187_
timestamp 1698431365
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1698431365
transform 1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1189_
timestamp 1698431365
transform 1 0 8096 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1698431365
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1191_
timestamp 1698431365
transform -1 0 8096 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1192_
timestamp 1698431365
transform -1 0 8740 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1698431365
transform 1 0 7636 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1194_
timestamp 1698431365
transform -1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1195_
timestamp 1698431365
transform -1 0 9476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1196_
timestamp 1698431365
transform 1 0 8188 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1197_
timestamp 1698431365
transform -1 0 8648 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 1698431365
transform 1 0 9476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1200_
timestamp 1698431365
transform -1 0 7176 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1698431365
transform 1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1202_
timestamp 1698431365
transform -1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1203_
timestamp 1698431365
transform -1 0 6256 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1698431365
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1205_
timestamp 1698431365
transform -1 0 7360 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1206_
timestamp 1698431365
transform -1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1207_
timestamp 1698431365
transform -1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1698431365
transform -1 0 9568 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1209_
timestamp 1698431365
transform 1 0 8004 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1698431365
transform 1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1698431365
transform 1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1698431365
transform 1 0 4600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1213_
timestamp 1698431365
transform -1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1698431365
transform 1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 1698431365
transform -1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1698431365
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1217_
timestamp 1698431365
transform 1 0 4232 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1218_
timestamp 1698431365
transform 1 0 4784 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1219_
timestamp 1698431365
transform 1 0 4324 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1220_
timestamp 1698431365
transform 1 0 4140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1221_
timestamp 1698431365
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1222_
timestamp 1698431365
transform -1 0 4968 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1698431365
transform -1 0 4876 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1224_
timestamp 1698431365
transform -1 0 3588 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1225_
timestamp 1698431365
transform -1 0 3220 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1698431365
transform 1 0 2300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1227_
timestamp 1698431365
transform 1 0 3036 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1698431365
transform 1 0 3220 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1229_
timestamp 1698431365
transform -1 0 4324 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1698431365
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1231_
timestamp 1698431365
transform -1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp 1698431365
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1233_
timestamp 1698431365
transform 1 0 3772 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1234_
timestamp 1698431365
transform 1 0 2760 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1235_
timestamp 1698431365
transform -1 0 2944 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1698431365
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1237_
timestamp 1698431365
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1238_
timestamp 1698431365
transform -1 0 8648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1239_
timestamp 1698431365
transform -1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1240_
timestamp 1698431365
transform -1 0 22540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1241_
timestamp 1698431365
transform -1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1698431365
transform -1 0 23920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 1698431365
transform -1 0 23552 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1244_
timestamp 1698431365
transform -1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1245_
timestamp 1698431365
transform 1 0 22632 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1246_
timestamp 1698431365
transform -1 0 23092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1247_
timestamp 1698431365
transform 1 0 23092 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1248_
timestamp 1698431365
transform -1 0 24288 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1249_
timestamp 1698431365
transform -1 0 24840 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1250_
timestamp 1698431365
transform 1 0 23552 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1698431365
transform 1 0 22540 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1698431365
transform 1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1253_
timestamp 1698431365
transform -1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1254_
timestamp 1698431365
transform 1 0 23368 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1255_
timestamp 1698431365
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1256_
timestamp 1698431365
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1257_
timestamp 1698431365
transform 1 0 24564 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1258_
timestamp 1698431365
transform -1 0 25208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1259_
timestamp 1698431365
transform -1 0 25300 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1260_
timestamp 1698431365
transform -1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1261_
timestamp 1698431365
transform -1 0 24288 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 24840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 1698431365
transform 1 0 5244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1698431365
transform 1 0 22724 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1265_
timestamp 1698431365
transform 1 0 21804 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1266_
timestamp 1698431365
transform -1 0 22724 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1267_
timestamp 1698431365
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1268_
timestamp 1698431365
transform -1 0 22724 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1698431365
transform -1 0 22632 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1270_
timestamp 1698431365
transform 1 0 21344 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1698431365
transform 1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1272_
timestamp 1698431365
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1698431365
transform 1 0 25392 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1274_
timestamp 1698431365
transform 1 0 24932 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1698431365
transform 1 0 26128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1276_
timestamp 1698431365
transform 1 0 23644 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1277_
timestamp 1698431365
transform -1 0 23276 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1278_
timestamp 1698431365
transform -1 0 24104 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1698431365
transform -1 0 23552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1280_
timestamp 1698431365
transform -1 0 24380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 1698431365
transform -1 0 21804 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11868 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 10580 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 1698431365
transform 1 0 12052 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1698431365
transform -1 0 11408 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 1698431365
transform 1 0 10212 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1698431365
transform -1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1288_
timestamp 1698431365
transform 1 0 19228 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1289_
timestamp 1698431365
transform 1 0 19136 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 1698431365
transform 1 0 17296 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1291_
timestamp 1698431365
transform 1 0 12052 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1292_
timestamp 1698431365
transform -1 0 16008 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1293_
timestamp 1698431365
transform -1 0 16008 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 14352 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1295_
timestamp 1698431365
transform 1 0 15456 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1296_
timestamp 1698431365
transform 1 0 17572 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1297_
timestamp 1698431365
transform 1 0 19228 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1298_
timestamp 1698431365
transform 1 0 19228 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1299_
timestamp 1698431365
transform 1 0 19320 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1300_
timestamp 1698431365
transform 1 0 19228 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 1698431365
transform 1 0 18768 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 1698431365
transform 1 0 14720 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1303_
timestamp 1698431365
transform 1 0 19044 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_2  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21804 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1306_
timestamp 1698431365
transform 1 0 16652 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1307_
timestamp 1698431365
transform 1 0 21620 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1308_
timestamp 1698431365
transform 1 0 21804 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1309_
timestamp 1698431365
transform -1 0 20608 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1310_
timestamp 1698431365
transform 1 0 19228 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1311_
timestamp 1698431365
transform -1 0 20056 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16652 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1313_
timestamp 1698431365
transform 1 0 13432 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1314_
timestamp 1698431365
transform -1 0 17848 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1315_
timestamp 1698431365
transform -1 0 17296 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1316_
timestamp 1698431365
transform 1 0 13340 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1317_
timestamp 1698431365
transform -1 0 11316 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 1698431365
transform 1 0 11316 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1319_
timestamp 1698431365
transform 1 0 2760 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1320_
timestamp 1698431365
transform -1 0 10488 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1321_
timestamp 1698431365
transform 1 0 4048 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1322_
timestamp 1698431365
transform 1 0 6900 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1323_
timestamp 1698431365
transform 1 0 6348 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1324_
timestamp 1698431365
transform 1 0 1380 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1325_
timestamp 1698431365
transform 1 0 1748 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1326_
timestamp 1698431365
transform 1 0 1472 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1327_
timestamp 1698431365
transform 1 0 6440 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1328_
timestamp 1698431365
transform 1 0 2300 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1329_
timestamp 1698431365
transform 1 0 6348 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 1698431365
transform 1 0 5888 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1331_
timestamp 1698431365
transform 1 0 1380 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1332_
timestamp 1698431365
transform 1 0 1564 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1333_
timestamp 1698431365
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1334_
timestamp 1698431365
transform 1 0 8096 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1335_
timestamp 1698431365
transform 1 0 3680 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1336_
timestamp 1698431365
transform 1 0 6716 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1698431365
transform 1 0 6348 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1338_
timestamp 1698431365
transform -1 0 3680 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1698431365
transform -1 0 4232 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1340_
timestamp 1698431365
transform 1 0 10120 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1341_
timestamp 1698431365
transform 1 0 9016 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1342_
timestamp 1698431365
transform 1 0 10028 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1343_
timestamp 1698431365
transform -1 0 16008 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1344_
timestamp 1698431365
transform -1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1345_
timestamp 1698431365
transform -1 0 18124 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 1698431365
transform 1 0 16652 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1347_
timestamp 1698431365
transform 1 0 19228 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1348_
timestamp 1698431365
transform 1 0 15824 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1349_
timestamp 1698431365
transform 1 0 18768 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1350_
timestamp 1698431365
transform 1 0 20608 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1351_
timestamp 1698431365
transform 1 0 19412 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1352_
timestamp 1698431365
transform -1 0 18584 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1353_
timestamp 1698431365
transform 1 0 14628 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1354_
timestamp 1698431365
transform 1 0 1564 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1355_
timestamp 1698431365
transform 1 0 9660 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1356_
timestamp 1698431365
transform 1 0 5152 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1357_
timestamp 1698431365
transform 1 0 9016 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 1698431365
transform 1 0 11592 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1359_
timestamp 1698431365
transform 1 0 1564 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1360_
timestamp 1698431365
transform 1 0 2300 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1698431365
transform -1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1698431365
transform 1 0 5796 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1698431365
transform 1 0 5152 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1698431365
transform 1 0 6256 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1698431365
transform 1 0 6532 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1366_
timestamp 1698431365
transform -1 0 16560 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1698431365
transform 1 0 1656 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1698431365
transform 1 0 1656 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1698431365
transform 1 0 3772 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1698431365
transform 1 0 1840 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1698431365
transform 1 0 1840 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1698431365
transform 1 0 8464 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1698431365
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1698431365
transform -1 0 23368 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1698431365
transform 1 0 24472 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1698431365
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1698431365
transform 1 0 24656 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1698431365
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1698431365
transform 1 0 20608 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1698431365
transform 1 0 21988 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1698431365
transform 1 0 24656 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1698431365
transform -1 0 24196 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1698431365
transform 1 0 24380 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1698431365
transform -1 0 22908 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK_SR $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14996 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform 1 0 13064 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLK_SR
timestamp 1698431365
transform -1 0 14812 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLK_SR
timestamp 1698431365
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform -1 0 9660 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform 1 0 16008 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform 1 0 18216 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform -1 0 7084 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform -1 0 7084 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform 1 0 15640 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_Dead_Time_Generator_inst_1.clk
timestamp 1698431365
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1698431365
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1698431365
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_63
timestamp 1698431365
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_75
timestamp 1698431365
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1698431365
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_94
timestamp 1698431365
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1698431365
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1698431365
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1698431365
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1698431365
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1698431365
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_147
timestamp 1698431365
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1698431365
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1698431365
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1698431365
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_181
timestamp 1698431365
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp 1698431365
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1698431365
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1698431365
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1698431365
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1698431365
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_225
timestamp 1698431365
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_232
timestamp 1698431365
transform 1 0 22448 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_244
timestamp 1698431365
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1698431365
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_265 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_275
timestamp 1698431365
transform 1 0 26404 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1698431365
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1698431365
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1698431365
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_71
timestamp 1698431365
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_76
timestamp 1698431365
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_82
timestamp 1698431365
transform 1 0 8648 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107
timestamp 1698431365
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1698431365
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1698431365
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1698431365
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_137
timestamp 1698431365
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_145
timestamp 1698431365
transform 1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_151
timestamp 1698431365
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_163
timestamp 1698431365
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1698431365
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_189
timestamp 1698431365
transform 1 0 18492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_201
timestamp 1698431365
transform 1 0 19596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_213
timestamp 1698431365
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 1698431365
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1698431365
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1698431365
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1698431365
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1698431365
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_273
timestamp 1698431365
transform 1 0 26220 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1698431365
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_15
timestamp 1698431365
transform 1 0 2484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_23
timestamp 1698431365
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_50
timestamp 1698431365
transform 1 0 5704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_59
timestamp 1698431365
transform 1 0 6532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_96
timestamp 1698431365
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_118
timestamp 1698431365
transform 1 0 11960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 1698431365
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_162
timestamp 1698431365
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_191
timestamp 1698431365
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1698431365
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1698431365
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1698431365
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1698431365
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1698431365
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1698431365
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1698431365
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1698431365
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1698431365
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1698431365
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1698431365
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_27
timestamp 1698431365
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_31
timestamp 1698431365
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_62
timestamp 1698431365
transform 1 0 6808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_74
timestamp 1698431365
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1698431365
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1698431365
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1698431365
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1698431365
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_216
timestamp 1698431365
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1698431365
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1698431365
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1698431365
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1698431365
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_273
timestamp 1698431365
transform 1 0 26220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1698431365
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1698431365
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1698431365
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1698431365
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_37
timestamp 1698431365
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_43
timestamp 1698431365
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_51
timestamp 1698431365
transform 1 0 5796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1698431365
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1698431365
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1698431365
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_119
timestamp 1698431365
transform 1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_123
timestamp 1698431365
transform 1 0 12420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_154
timestamp 1698431365
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_161
timestamp 1698431365
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_179
timestamp 1698431365
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_183
timestamp 1698431365
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1698431365
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_218
timestamp 1698431365
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_230
timestamp 1698431365
transform 1 0 22264 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_242
timestamp 1698431365
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1698431365
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1698431365
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1698431365
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1698431365
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_17
timestamp 1698431365
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_29
timestamp 1698431365
transform 1 0 3772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_41
timestamp 1698431365
transform 1 0 4876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_49
timestamp 1698431365
transform 1 0 5612 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1698431365
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_69
timestamp 1698431365
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1698431365
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1698431365
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1698431365
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 1698431365
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_121
timestamp 1698431365
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_126
timestamp 1698431365
transform 1 0 12696 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_155
timestamp 1698431365
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1698431365
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1698431365
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1698431365
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_193
timestamp 1698431365
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_200
timestamp 1698431365
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_207
timestamp 1698431365
transform 1 0 20148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_219
timestamp 1698431365
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1698431365
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1698431365
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1698431365
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1698431365
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1698431365
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_273
timestamp 1698431365
transform 1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1698431365
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1698431365
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1698431365
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1698431365
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_41
timestamp 1698431365
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_50
timestamp 1698431365
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_60
timestamp 1698431365
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_72
timestamp 1698431365
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1698431365
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1698431365
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1698431365
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1698431365
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1698431365
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_182
timestamp 1698431365
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1698431365
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 1698431365
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_205
timestamp 1698431365
transform 1 0 19964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_217
timestamp 1698431365
transform 1 0 21068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_229
timestamp 1698431365
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_241
timestamp 1698431365
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1698431365
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1698431365
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_265
timestamp 1698431365
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_269
timestamp 1698431365
transform 1 0 25852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_6
timestamp 1698431365
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_34
timestamp 1698431365
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_86
timestamp 1698431365
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1698431365
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1698431365
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1698431365
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1698431365
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_149
timestamp 1698431365
transform 1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_154
timestamp 1698431365
transform 1 0 15272 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_162
timestamp 1698431365
transform 1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1698431365
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1698431365
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_174
timestamp 1698431365
transform 1 0 17112 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_186
timestamp 1698431365
transform 1 0 18216 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_194
timestamp 1698431365
transform 1 0 18952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_205
timestamp 1698431365
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_211
timestamp 1698431365
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1698431365
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_228
timestamp 1698431365
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_240
timestamp 1698431365
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_252
timestamp 1698431365
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_264
timestamp 1698431365
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_276
timestamp 1698431365
transform 1 0 26496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1698431365
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1698431365
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_69
timestamp 1698431365
transform 1 0 7452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_75
timestamp 1698431365
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1698431365
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_92
timestamp 1698431365
transform 1 0 9568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_125
timestamp 1698431365
transform 1 0 12604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1698431365
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1698431365
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_153
timestamp 1698431365
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_159
timestamp 1698431365
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_189
timestamp 1698431365
transform 1 0 18492 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1698431365
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1698431365
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1698431365
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1698431365
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1698431365
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1698431365
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1698431365
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_19
timestamp 1698431365
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_29
timestamp 1698431365
transform 1 0 3772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1698431365
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1698431365
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 1698431365
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_125
timestamp 1698431365
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1698431365
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1698431365
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1698431365
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1698431365
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_183
timestamp 1698431365
transform 1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1698431365
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1698431365
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1698431365
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1698431365
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_273
timestamp 1698431365
transform 1 0 26220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1698431365
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_14
timestamp 1698431365
transform 1 0 2392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1698431365
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1698431365
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_65
timestamp 1698431365
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_69
timestamp 1698431365
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1698431365
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1698431365
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_90
timestamp 1698431365
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_102
timestamp 1698431365
transform 1 0 10488 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_115
timestamp 1698431365
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_132
timestamp 1698431365
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_144
timestamp 1698431365
transform 1 0 14352 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_161
timestamp 1698431365
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_173
timestamp 1698431365
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1698431365
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_216
timestamp 1698431365
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_228
timestamp 1698431365
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_240
timestamp 1698431365
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1698431365
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1698431365
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1698431365
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1698431365
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1698431365
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1698431365
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1698431365
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1698431365
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1698431365
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1698431365
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_86
timestamp 1698431365
transform 1 0 9016 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_98
timestamp 1698431365
transform 1 0 10120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1698431365
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1698431365
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_125
timestamp 1698431365
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_147
timestamp 1698431365
transform 1 0 14628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_159
timestamp 1698431365
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1698431365
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1698431365
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 1698431365
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_198
timestamp 1698431365
transform 1 0 19320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_225
timestamp 1698431365
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_231
timestamp 1698431365
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_251
timestamp 1698431365
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_263
timestamp 1698431365
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_275
timestamp 1698431365
transform 1 0 26404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_6
timestamp 1698431365
transform 1 0 1656 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_20
timestamp 1698431365
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_36
timestamp 1698431365
transform 1 0 4416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_48
timestamp 1698431365
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_55
timestamp 1698431365
transform 1 0 6164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_67
timestamp 1698431365
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_74
timestamp 1698431365
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1698431365
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1698431365
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_97
timestamp 1698431365
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_110
timestamp 1698431365
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_137
timestamp 1698431365
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1698431365
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_153
timestamp 1698431365
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_160
timestamp 1698431365
transform 1 0 15824 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_200
timestamp 1698431365
transform 1 0 19504 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_208
timestamp 1698431365
transform 1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_213
timestamp 1698431365
transform 1 0 20700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_219
timestamp 1698431365
transform 1 0 21252 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1698431365
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1698431365
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_265
timestamp 1698431365
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_269
timestamp 1698431365
transform 1 0 25852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1698431365
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 1698431365
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_41
timestamp 1698431365
transform 1 0 4876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_49
timestamp 1698431365
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_69
timestamp 1698431365
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_85
timestamp 1698431365
transform 1 0 8924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_97
timestamp 1698431365
transform 1 0 10028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_101
timestamp 1698431365
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1698431365
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_116
timestamp 1698431365
transform 1 0 11776 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_128
timestamp 1698431365
transform 1 0 12880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_140
timestamp 1698431365
transform 1 0 13984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_146
timestamp 1698431365
transform 1 0 14536 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_190
timestamp 1698431365
transform 1 0 18584 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_202
timestamp 1698431365
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_214
timestamp 1698431365
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_218
timestamp 1698431365
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1698431365
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_244
timestamp 1698431365
transform 1 0 23552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_250
timestamp 1698431365
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_258
timestamp 1698431365
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_269
timestamp 1698431365
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1698431365
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1698431365
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1698431365
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1698431365
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_91
timestamp 1698431365
transform 1 0 9476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1698431365
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_148
timestamp 1698431365
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_160
timestamp 1698431365
transform 1 0 15824 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_172
timestamp 1698431365
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_184
timestamp 1698431365
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1698431365
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_209
timestamp 1698431365
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1698431365
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_275
timestamp 1698431365
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1698431365
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_50
timestamp 1698431365
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_60
timestamp 1698431365
transform 1 0 6624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_83
timestamp 1698431365
transform 1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_121
timestamp 1698431365
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_129
timestamp 1698431365
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_137
timestamp 1698431365
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_141
timestamp 1698431365
transform 1 0 14076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_157
timestamp 1698431365
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1698431365
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1698431365
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1698431365
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_193
timestamp 1698431365
transform 1 0 18860 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_199
timestamp 1698431365
transform 1 0 19412 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_203
timestamp 1698431365
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_215
timestamp 1698431365
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1698431365
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_238
timestamp 1698431365
transform 1 0 23000 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_246
timestamp 1698431365
transform 1 0 23736 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_269
timestamp 1698431365
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1698431365
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1698431365
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1698431365
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_41
timestamp 1698431365
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1698431365
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1698431365
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1698431365
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1698431365
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp 1698431365
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_99
timestamp 1698431365
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1698431365
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_188
timestamp 1698431365
transform 1 0 18400 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_192
timestamp 1698431365
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_220
timestamp 1698431365
transform 1 0 21344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_229
timestamp 1698431365
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_238
timestamp 1698431365
transform 1 0 23000 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1698431365
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1698431365
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_257
timestamp 1698431365
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_266
timestamp 1698431365
transform 1 0 25576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_274
timestamp 1698431365
transform 1 0 26312 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1698431365
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1698431365
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1698431365
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1698431365
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1698431365
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1698431365
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1698431365
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1698431365
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1698431365
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1698431365
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1698431365
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1698431365
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1698431365
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_125
timestamp 1698431365
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_132
timestamp 1698431365
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_172
timestamp 1698431365
transform 1 0 16928 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_202
timestamp 1698431365
transform 1 0 19688 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_208
timestamp 1698431365
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1698431365
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_225
timestamp 1698431365
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_250
timestamp 1698431365
transform 1 0 24104 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_263
timestamp 1698431365
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_271
timestamp 1698431365
transform 1 0 26036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1698431365
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1698431365
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_20
timestamp 1698431365
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_40
timestamp 1698431365
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_52
timestamp 1698431365
transform 1 0 5888 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_64
timestamp 1698431365
transform 1 0 6992 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_76
timestamp 1698431365
transform 1 0 8096 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1698431365
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1698431365
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1698431365
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_109
timestamp 1698431365
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_114
timestamp 1698431365
transform 1 0 11592 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1698431365
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1698431365
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_153
timestamp 1698431365
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_176
timestamp 1698431365
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_188
timestamp 1698431365
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1698431365
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_220
timestamp 1698431365
transform 1 0 21344 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_227
timestamp 1698431365
transform 1 0 21988 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_233
timestamp 1698431365
transform 1 0 22540 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_240
timestamp 1698431365
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1698431365
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1698431365
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1698431365
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1698431365
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_33
timestamp 1698431365
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_49
timestamp 1698431365
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1698431365
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1698431365
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 1698431365
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_90
timestamp 1698431365
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_122
timestamp 1698431365
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 1698431365
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 1698431365
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_169
timestamp 1698431365
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_177
timestamp 1698431365
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_198
timestamp 1698431365
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_213
timestamp 1698431365
transform 1 0 20700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1698431365
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_228
timestamp 1698431365
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_240
timestamp 1698431365
transform 1 0 23184 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_266
timestamp 1698431365
transform 1 0 25576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_276
timestamp 1698431365
transform 1 0 26496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1698431365
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_24
timestamp 1698431365
transform 1 0 3312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_49
timestamp 1698431365
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_67
timestamp 1698431365
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_132
timestamp 1698431365
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1698431365
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_154
timestamp 1698431365
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_166
timestamp 1698431365
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_178
timestamp 1698431365
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_182
timestamp 1698431365
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_188
timestamp 1698431365
transform 1 0 18400 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_197
timestamp 1698431365
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1698431365
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_233
timestamp 1698431365
transform 1 0 22540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_241
timestamp 1698431365
transform 1 0 23276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_253
timestamp 1698431365
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_272
timestamp 1698431365
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_276
timestamp 1698431365
transform 1 0 26496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_6
timestamp 1698431365
transform 1 0 1656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2208 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_20
timestamp 1698431365
transform 1 0 2944 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_32
timestamp 1698431365
transform 1 0 4048 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_39
timestamp 1698431365
transform 1 0 4692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1698431365
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1698431365
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_74
timestamp 1698431365
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_83
timestamp 1698431365
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_98
timestamp 1698431365
transform 1 0 10120 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_104
timestamp 1698431365
transform 1 0 10672 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 1698431365
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_116
timestamp 1698431365
transform 1 0 11776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_158
timestamp 1698431365
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1698431365
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_169
timestamp 1698431365
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_180
timestamp 1698431365
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_184
timestamp 1698431365
transform 1 0 18032 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_191
timestamp 1698431365
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_203
timestamp 1698431365
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_215
timestamp 1698431365
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1698431365
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_225
timestamp 1698431365
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 23552 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_257
timestamp 1698431365
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_263
timestamp 1698431365
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_267
timestamp 1698431365
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_276
timestamp 1698431365
transform 1 0 26496 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1698431365
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_15
timestamp 1698431365
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1698431365
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1698431365
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_53
timestamp 1698431365
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_61
timestamp 1698431365
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_66
timestamp 1698431365
transform 1 0 7176 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_76
timestamp 1698431365
transform 1 0 8096 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1698431365
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_94
timestamp 1698431365
transform 1 0 9752 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_106
timestamp 1698431365
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_118
timestamp 1698431365
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_131
timestamp 1698431365
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1698431365
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_156
timestamp 1698431365
transform 1 0 15456 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_162
timestamp 1698431365
transform 1 0 16008 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_200
timestamp 1698431365
transform 1 0 19504 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_208
timestamp 1698431365
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_220
timestamp 1698431365
transform 1 0 21344 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_228
timestamp 1698431365
transform 1 0 22080 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 23552 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1698431365
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_271
timestamp 1698431365
transform 1 0 26036 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1698431365
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_15
timestamp 1698431365
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_26
timestamp 1698431365
transform 1 0 3496 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_38
timestamp 1698431365
transform 1 0 4600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_46
timestamp 1698431365
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1698431365
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1698431365
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1698431365
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1698431365
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1698431365
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1698431365
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1698431365
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_125
timestamp 1698431365
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1698431365
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_150
timestamp 1698431365
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1698431365
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_172
timestamp 1698431365
transform 1 0 16928 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_196
timestamp 1698431365
transform 1 0 19136 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_218
timestamp 1698431365
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1698431365
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_233
timestamp 1698431365
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_237
timestamp 1698431365
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_241
timestamp 1698431365
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_247
timestamp 1698431365
transform 1 0 23828 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_262
timestamp 1698431365
transform 1 0 25208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_276
timestamp 1698431365
transform 1 0 26496 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_6
timestamp 1698431365
transform 1 0 1656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_12
timestamp 1698431365
transform 1 0 2208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_41
timestamp 1698431365
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_75
timestamp 1698431365
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1698431365
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1698431365
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_97
timestamp 1698431365
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_119
timestamp 1698431365
transform 1 0 12052 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_128
timestamp 1698431365
transform 1 0 12880 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_132
timestamp 1698431365
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1698431365
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_149
timestamp 1698431365
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_183
timestamp 1698431365
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1698431365
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_205
timestamp 1698431365
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_217
timestamp 1698431365
transform 1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_224
timestamp 1698431365
transform 1 0 21712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1698431365
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_253
timestamp 1698431365
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_270
timestamp 1698431365
transform 1 0 25944 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_276
timestamp 1698431365
transform 1 0 26496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_22
timestamp 1698431365
transform 1 0 3128 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_43
timestamp 1698431365
transform 1 0 5060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 1698431365
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1698431365
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_78
timestamp 1698431365
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_102
timestamp 1698431365
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_117
timestamp 1698431365
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_177
timestamp 1698431365
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_187
timestamp 1698431365
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_192
timestamp 1698431365
transform 1 0 18768 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_253
timestamp 1698431365
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_262
timestamp 1698431365
transform 1 0 25208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_274
timestamp 1698431365
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_3
timestamp 1698431365
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1698431365
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_48
timestamp 1698431365
transform 1 0 5520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_72
timestamp 1698431365
transform 1 0 7728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_96
timestamp 1698431365
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_115
timestamp 1698431365
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1698431365
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1698431365
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_149
timestamp 1698431365
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_183
timestamp 1698431365
transform 1 0 17940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1698431365
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_204
timestamp 1698431365
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_211
timestamp 1698431365
transform 1 0 20516 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_219
timestamp 1698431365
transform 1 0 21252 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_238
timestamp 1698431365
transform 1 0 23000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1698431365
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1698431365
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1698431365
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1698431365
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1698431365
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_27
timestamp 1698431365
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_34
timestamp 1698431365
transform 1 0 4232 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1698431365
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_81
timestamp 1698431365
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1698431365
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_116
timestamp 1698431365
transform 1 0 11776 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_148
timestamp 1698431365
transform 1 0 14720 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_152
timestamp 1698431365
transform 1 0 15088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_162
timestamp 1698431365
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_172
timestamp 1698431365
transform 1 0 16928 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_184
timestamp 1698431365
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1698431365
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1698431365
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1698431365
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_233
timestamp 1698431365
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_239
timestamp 1698431365
transform 1 0 23092 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_251
timestamp 1698431365
transform 1 0 24196 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_263
timestamp 1698431365
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_275
timestamp 1698431365
transform 1 0 26404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_6
timestamp 1698431365
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_18
timestamp 1698431365
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1698431365
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1698431365
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_41
timestamp 1698431365
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1698431365
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1698431365
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1698431365
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1698431365
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1698431365
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1698431365
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_121
timestamp 1698431365
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_127
timestamp 1698431365
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_131
timestamp 1698431365
transform 1 0 13156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1698431365
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_157
timestamp 1698431365
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_178
timestamp 1698431365
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_186
timestamp 1698431365
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1698431365
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1698431365
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1698431365
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_237
timestamp 1698431365
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1698431365
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1698431365
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1698431365
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1698431365
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_11
timestamp 1698431365
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_34
timestamp 1698431365
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_46
timestamp 1698431365
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1698431365
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1698431365
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1698431365
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1698431365
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_93
timestamp 1698431365
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_98
timestamp 1698431365
transform 1 0 10120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1698431365
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1698431365
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_125
timestamp 1698431365
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_153
timestamp 1698431365
transform 1 0 15180 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1698431365
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_180
timestamp 1698431365
transform 1 0 17664 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_192
timestamp 1698431365
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_203
timestamp 1698431365
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 1698431365
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1698431365
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1698431365
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1698431365
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1698431365
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1698431365
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_273
timestamp 1698431365
transform 1 0 26220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1698431365
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1698431365
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_36
timestamp 1698431365
transform 1 0 4416 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_47
timestamp 1698431365
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_59
timestamp 1698431365
transform 1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1698431365
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1698431365
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1698431365
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_98
timestamp 1698431365
transform 1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_108
timestamp 1698431365
transform 1 0 11040 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_120
timestamp 1698431365
transform 1 0 12144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_129
timestamp 1698431365
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1698431365
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_165
timestamp 1698431365
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1698431365
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_212
timestamp 1698431365
transform 1 0 20608 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_224
timestamp 1698431365
transform 1 0 21712 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_236
timestamp 1698431365
transform 1 0 22816 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_248
timestamp 1698431365
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1698431365
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_265
timestamp 1698431365
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 1698431365
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_11
timestamp 1698431365
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_17
timestamp 1698431365
transform 1 0 2668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_22
timestamp 1698431365
transform 1 0 3128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_30
timestamp 1698431365
transform 1 0 3864 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1698431365
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_80
timestamp 1698431365
transform 1 0 8464 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1698431365
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1698431365
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_121
timestamp 1698431365
transform 1 0 12236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_133
timestamp 1698431365
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_140
timestamp 1698431365
transform 1 0 13984 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_149
timestamp 1698431365
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_153
timestamp 1698431365
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_174
timestamp 1698431365
transform 1 0 17112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1698431365
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1698431365
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1698431365
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1698431365
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1698431365
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1698431365
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_273
timestamp 1698431365
transform 1 0 26220 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1698431365
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_18
timestamp 1698431365
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1698431365
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1698431365
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_37
timestamp 1698431365
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_43
timestamp 1698431365
transform 1 0 5060 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_49
timestamp 1698431365
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_61
timestamp 1698431365
transform 1 0 6716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_65
timestamp 1698431365
transform 1 0 7084 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_69
timestamp 1698431365
transform 1 0 7452 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_77
timestamp 1698431365
transform 1 0 8188 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1698431365
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_93
timestamp 1698431365
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 10672 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_122
timestamp 1698431365
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_129
timestamp 1698431365
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1698431365
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 1698431365
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_168
timestamp 1698431365
transform 1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_189
timestamp 1698431365
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_218
timestamp 1698431365
transform 1 0 21160 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_230
timestamp 1698431365
transform 1 0 22264 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_242
timestamp 1698431365
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1698431365
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1698431365
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1698431365
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1698431365
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_15
timestamp 1698431365
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp 1698431365
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_33
timestamp 1698431365
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1698431365
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1698431365
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_108
timestamp 1698431365
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_118
timestamp 1698431365
transform 1 0 11960 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_130
timestamp 1698431365
transform 1 0 13064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_142
timestamp 1698431365
transform 1 0 14168 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_150
timestamp 1698431365
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1698431365
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_197
timestamp 1698431365
transform 1 0 19228 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_203
timestamp 1698431365
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_207
timestamp 1698431365
transform 1 0 20148 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_219
timestamp 1698431365
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1698431365
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1698431365
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1698431365
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1698431365
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1698431365
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_273
timestamp 1698431365
transform 1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_3
timestamp 1698431365
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 1698431365
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1698431365
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1698431365
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1698431365
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1698431365
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_89
timestamp 1698431365
transform 1 0 9292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_93
timestamp 1698431365
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_102
timestamp 1698431365
transform 1 0 10488 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_114
timestamp 1698431365
transform 1 0 11592 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_126
timestamp 1698431365
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_131
timestamp 1698431365
transform 1 0 13156 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_150
timestamp 1698431365
transform 1 0 14904 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_181
timestamp 1698431365
transform 1 0 17756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1698431365
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1698431365
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1698431365
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1698431365
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1698431365
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1698431365
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1698431365
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1698431365
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1698431365
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_41
timestamp 1698431365
transform 1 0 4876 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_67
timestamp 1698431365
transform 1 0 7268 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_79
timestamp 1698431365
transform 1 0 8372 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_91
timestamp 1698431365
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_103
timestamp 1698431365
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1698431365
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1698431365
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1698431365
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1698431365
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1698431365
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_187
timestamp 1698431365
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_199
timestamp 1698431365
transform 1 0 19412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_211
timestamp 1698431365
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1698431365
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1698431365
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1698431365
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1698431365
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1698431365
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_273
timestamp 1698431365
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_6
timestamp 1698431365
transform 1 0 1656 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1698431365
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_47
timestamp 1698431365
transform 1 0 5428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_51
timestamp 1698431365
transform 1 0 5796 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_72
timestamp 1698431365
transform 1 0 7728 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_93
timestamp 1698431365
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_99
timestamp 1698431365
transform 1 0 10212 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_107
timestamp 1698431365
transform 1 0 10948 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_122
timestamp 1698431365
transform 1 0 12328 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_134
timestamp 1698431365
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_162
timestamp 1698431365
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_169
timestamp 1698431365
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_173
timestamp 1698431365
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_177
timestamp 1698431365
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_186
timestamp 1698431365
transform 1 0 18216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1698431365
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_207
timestamp 1698431365
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_216
timestamp 1698431365
transform 1 0 20976 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_226
timestamp 1698431365
transform 1 0 21896 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_232
timestamp 1698431365
transform 1 0 22448 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_236
timestamp 1698431365
transform 1 0 22816 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 1698431365
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1698431365
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1698431365
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1698431365
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1698431365
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1698431365
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1698431365
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1698431365
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1698431365
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1698431365
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_69
timestamp 1698431365
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_77
timestamp 1698431365
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_99
timestamp 1698431365
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1698431365
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_129
timestamp 1698431365
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_155
timestamp 1698431365
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_159
timestamp 1698431365
transform 1 0 15732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1698431365
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1698431365
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_248
timestamp 1698431365
transform 1 0 23920 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_260
timestamp 1698431365
transform 1 0 25024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_272
timestamp 1698431365
transform 1 0 26128 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_276
timestamp 1698431365
transform 1 0 26496 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1698431365
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_15
timestamp 1698431365
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_24
timestamp 1698431365
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1698431365
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_41
timestamp 1698431365
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_49
timestamp 1698431365
transform 1 0 5612 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_57
timestamp 1698431365
transform 1 0 6348 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_63
timestamp 1698431365
transform 1 0 6900 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_67
timestamp 1698431365
transform 1 0 7268 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_75
timestamp 1698431365
transform 1 0 8004 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_120
timestamp 1698431365
transform 1 0 12144 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1698431365
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1698431365
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_153
timestamp 1698431365
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_176
timestamp 1698431365
transform 1 0 17296 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_184
timestamp 1698431365
transform 1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_209
timestamp 1698431365
transform 1 0 20332 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1698431365
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1698431365
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1698431365
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_6
timestamp 1698431365
transform 1 0 1656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2024 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_20
timestamp 1698431365
transform 1 0 2944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_28
timestamp 1698431365
transform 1 0 3680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_34
timestamp 1698431365
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_46
timestamp 1698431365
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1698431365
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_78
timestamp 1698431365
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_86
timestamp 1698431365
transform 1 0 9016 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1698431365
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_125
timestamp 1698431365
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_133
timestamp 1698431365
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_140
timestamp 1698431365
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_155
timestamp 1698431365
transform 1 0 15364 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_163
timestamp 1698431365
transform 1 0 16100 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1698431365
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1698431365
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1698431365
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_193
timestamp 1698431365
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1698431365
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_217
timestamp 1698431365
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1698431365
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1698431365
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1698431365
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_273
timestamp 1698431365
transform 1 0 26220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1698431365
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_29
timestamp 1698431365
transform 1 0 3772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_45
timestamp 1698431365
transform 1 0 5244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_53
timestamp 1698431365
transform 1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_68
timestamp 1698431365
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1698431365
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1698431365
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_101
timestamp 1698431365
transform 1 0 10396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_113
timestamp 1698431365
transform 1 0 11500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_125
timestamp 1698431365
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1698431365
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1698431365
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1698431365
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1698431365
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1698431365
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1698431365
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1698431365
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_207
timestamp 1698431365
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_219
timestamp 1698431365
transform 1 0 21252 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_223
timestamp 1698431365
transform 1 0 21620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_232
timestamp 1698431365
transform 1 0 22448 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_242
timestamp 1698431365
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1698431365
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1698431365
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1698431365
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1698431365
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_51
timestamp 1698431365
transform 1 0 5796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_64
timestamp 1698431365
transform 1 0 6992 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_79
timestamp 1698431365
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_91
timestamp 1698431365
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_103
timestamp 1698431365
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1698431365
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1698431365
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_140
timestamp 1698431365
transform 1 0 13984 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_148
timestamp 1698431365
transform 1 0 14720 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_158
timestamp 1698431365
transform 1 0 15640 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_164
timestamp 1698431365
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1698431365
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_181
timestamp 1698431365
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_212
timestamp 1698431365
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_246
timestamp 1698431365
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_258
timestamp 1698431365
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_270
timestamp 1698431365
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_276
timestamp 1698431365
transform 1 0 26496 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1698431365
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1698431365
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1698431365
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_44
timestamp 1698431365
transform 1 0 5152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_56
timestamp 1698431365
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_68
timestamp 1698431365
transform 1 0 7360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1698431365
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1698431365
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_105
timestamp 1698431365
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_128
timestamp 1698431365
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_132
timestamp 1698431365
transform 1 0 13248 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_148
timestamp 1698431365
transform 1 0 14720 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_171
timestamp 1698431365
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_183
timestamp 1698431365
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1698431365
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_204
timestamp 1698431365
transform 1 0 19872 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_216
timestamp 1698431365
transform 1 0 20976 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_228
timestamp 1698431365
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_240
timestamp 1698431365
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1698431365
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1698431365
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1698431365
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_15
timestamp 1698431365
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_45
timestamp 1698431365
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_53
timestamp 1698431365
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_57
timestamp 1698431365
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_75
timestamp 1698431365
transform 1 0 8004 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_102
timestamp 1698431365
transform 1 0 10488 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_113
timestamp 1698431365
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_154
timestamp 1698431365
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_158
timestamp 1698431365
transform 1 0 15640 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1698431365
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_190
timestamp 1698431365
transform 1 0 18584 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_198
timestamp 1698431365
transform 1 0 19320 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_203
timestamp 1698431365
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_215
timestamp 1698431365
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1698431365
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1698431365
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1698431365
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1698431365
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1698431365
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_273
timestamp 1698431365
transform 1 0 26220 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1698431365
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_15
timestamp 1698431365
transform 1 0 2484 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_23
timestamp 1698431365
transform 1 0 3220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_53
timestamp 1698431365
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_88
timestamp 1698431365
transform 1 0 9200 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_131
timestamp 1698431365
transform 1 0 13156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_150
timestamp 1698431365
transform 1 0 14904 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_156
timestamp 1698431365
transform 1 0 15456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_185
timestamp 1698431365
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_220
timestamp 1698431365
transform 1 0 21344 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_232
timestamp 1698431365
transform 1 0 22448 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_244
timestamp 1698431365
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1698431365
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1698431365
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1698431365
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_27
timestamp 1698431365
transform 1 0 3588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_45
timestamp 1698431365
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_53
timestamp 1698431365
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_57
timestamp 1698431365
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_71
timestamp 1698431365
transform 1 0 7636 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_83
timestamp 1698431365
transform 1 0 8740 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_95
timestamp 1698431365
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_102
timestamp 1698431365
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_106
timestamp 1698431365
transform 1 0 10856 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1698431365
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1698431365
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_128
timestamp 1698431365
transform 1 0 12880 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_132
timestamp 1698431365
transform 1 0 13248 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_144
timestamp 1698431365
transform 1 0 14352 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_156
timestamp 1698431365
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_180
timestamp 1698431365
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_184
timestamp 1698431365
transform 1 0 18032 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_206
timestamp 1698431365
transform 1 0 20056 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_218
timestamp 1698431365
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1698431365
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1698431365
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1698431365
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1698431365
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_273
timestamp 1698431365
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1698431365
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1698431365
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1698431365
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_35
timestamp 1698431365
transform 1 0 4324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_47
timestamp 1698431365
transform 1 0 5428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_55
timestamp 1698431365
transform 1 0 6164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_57
timestamp 1698431365
transform 1 0 6348 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_66
timestamp 1698431365
transform 1 0 7176 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_78
timestamp 1698431365
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1698431365
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_97
timestamp 1698431365
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_101
timestamp 1698431365
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_108
timestamp 1698431365
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1698431365
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 1698431365
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1698431365
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1698431365
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1698431365
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1698431365
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_169
timestamp 1698431365
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_177
timestamp 1698431365
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_184
timestamp 1698431365
transform 1 0 18032 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1698431365
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1698431365
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 1698431365
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1698431365
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1698431365
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1698431365
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_253
timestamp 1698431365
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_260
timestamp 1698431365
transform 1 0 25024 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_272
timestamp 1698431365
transform 1 0 26128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_276
timestamp 1698431365
transform 1 0 26496 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  hold2
timestamp 1698431365
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 24748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1698431365
transform -1 0 24104 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1698431365
transform -1 0 25576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1698431365
transform 1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1698431365
transform -1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1698431365
transform -1 0 26496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1698431365
transform -1 0 9936 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1698431365
transform -1 0 9108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1698431365
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1698431365
transform -1 0 23828 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1698431365
transform 1 0 21804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1698431365
transform -1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1698431365
transform -1 0 8280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1698431365
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1698431365
transform -1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1698431365
transform -1 0 15364 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1698431365
transform 1 0 9108 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1698431365
transform 1 0 25760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1698431365
transform -1 0 11316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1698431365
transform -1 0 18492 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1698431365
transform -1 0 21712 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1698431365
transform -1 0 7912 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1698431365
transform 1 0 23276 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold26
timestamp 1698431365
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  hold27
timestamp 1698431365
transform -1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1698431365
transform 1 0 12604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17388 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1698431365
transform -1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1698431365
transform 1 0 9016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1698431365
transform -1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1698431365
transform -1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1698431365
transform -1 0 5796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1698431365
transform -1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1698431365
transform 1 0 4232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1698431365
transform -1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1698431365
transform -1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1698431365
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1698431365
transform 1 0 3864 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1698431365
transform -1 0 5060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1698431365
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1698431365
transform -1 0 19964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1698431365
transform 1 0 5796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1698431365
transform -1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1698431365
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1698431365
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1698431365
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1698431365
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1698431365
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1698431365
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1698431365
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1698431365
transform 1 0 26312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1698431365
transform -1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1698431365
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1698431365
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1698431365
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1698431365
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1698431365
transform 1 0 24472 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1698431365
transform 1 0 17940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1698431365
transform -1 0 11040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1698431365
transform -1 0 10580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1698431365
transform 1 0 25852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1698431365
transform -1 0 4324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1698431365
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1698431365
transform 1 0 17480 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1698431365
transform -1 0 14628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1698431365
transform 1 0 21896 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  output25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1698431365
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1698431365
transform -1 0 26864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1698431365
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1698431365
transform -1 0 26864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1698431365
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1698431365
transform -1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1698431365
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1698431365
transform -1 0 26864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1698431365
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1698431365
transform -1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1698431365
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1698431365
transform -1 0 26864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1698431365
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1698431365
transform -1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1698431365
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1698431365
transform -1 0 26864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1698431365
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1698431365
transform -1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1698431365
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1698431365
transform -1 0 26864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1698431365
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1698431365
transform -1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1698431365
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1698431365
transform -1 0 26864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1698431365
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1698431365
transform -1 0 26864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1698431365
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1698431365
transform -1 0 26864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1698431365
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1698431365
transform -1 0 26864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1698431365
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1698431365
transform -1 0 26864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1698431365
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1698431365
transform -1 0 26864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1698431365
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1698431365
transform -1 0 26864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1698431365
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1698431365
transform -1 0 26864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1698431365
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1698431365
transform -1 0 26864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1698431365
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1698431365
transform -1 0 26864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1698431365
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1698431365
transform -1 0 26864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1698431365
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1698431365
transform -1 0 26864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1698431365
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1698431365
transform -1 0 26864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1698431365
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1698431365
transform -1 0 26864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1698431365
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1698431365
transform -1 0 26864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1698431365
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1698431365
transform -1 0 26864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1698431365
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1698431365
transform -1 0 26864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1698431365
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1698431365
transform -1 0 26864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1698431365
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1698431365
transform -1 0 26864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1698431365
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1698431365
transform -1 0 26864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1698431365
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1698431365
transform -1 0 26864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1698431365
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1698431365
transform -1 0 26864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1698431365
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1698431365
transform -1 0 26864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1698431365
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1698431365
transform -1 0 26864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1698431365
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1698431365
transform -1 0 26864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1698431365
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1698431365
transform -1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1698431365
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1698431365
transform -1 0 26864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1698431365
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1698431365
transform -1 0 26864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1698431365
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1698431365
transform -1 0 26864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1698431365
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1698431365
transform -1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1698431365
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1698431365
transform -1 0 26864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1698431365
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1698431365
transform -1 0 26864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1698431365
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1698431365
transform -1 0 26864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1698431365
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1698431365
transform -1 0 26864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1698431365
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1698431365
transform -1 0 26864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1698431365
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1698431365
transform -1 0 26864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  rebuffer1
timestamp 1698431365
transform 1 0 14168 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1698431365
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1698431365
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1698431365
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1698431365
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1698431365
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1698431365
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1698431365
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1698431365
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1698431365
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1698431365
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1698431365
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1698431365
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1698431365
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1698431365
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1698431365
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1698431365
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1698431365
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1698431365
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1698431365
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1698431365
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1698431365
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1698431365
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1698431365
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1698431365
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1698431365
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1698431365
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1698431365
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1698431365
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1698431365
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1698431365
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1698431365
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1698431365
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1698431365
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1698431365
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1698431365
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1698431365
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1698431365
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1698431365
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1698431365
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1698431365
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1698431365
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1698431365
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1698431365
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1698431365
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1698431365
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1698431365
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1698431365
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1698431365
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1698431365
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1698431365
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1698431365
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1698431365
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1698431365
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1698431365
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1698431365
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1698431365
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1698431365
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1698431365
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1698431365
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1698431365
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1698431365
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1698431365
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1698431365
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1698431365
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1698431365
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1698431365
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1698431365
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1698431365
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1698431365
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1698431365
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1698431365
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1698431365
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1698431365
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1698431365
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1698431365
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1698431365
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1698431365
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1698431365
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1698431365
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1698431365
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1698431365
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1698431365
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1698431365
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1698431365
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1698431365
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1698431365
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1698431365
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1698431365
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1698431365
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1698431365
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1698431365
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1698431365
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1698431365
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1698431365
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1698431365
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1698431365
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1698431365
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1698431365
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1698431365
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1698431365
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1698431365
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1698431365
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1698431365
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1698431365
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1698431365
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1698431365
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1698431365
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1698431365
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1698431365
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1698431365
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1698431365
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1698431365
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1698431365
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1698431365
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1698431365
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1698431365
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1698431365
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1698431365
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1698431365
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1698431365
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1698431365
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1698431365
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1698431365
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1698431365
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1698431365
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1698431365
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1698431365
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1698431365
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1698431365
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1698431365
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1698431365
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1698431365
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1698431365
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1698431365
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1698431365
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1698431365
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1698431365
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1698431365
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1698431365
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1698431365
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1698431365
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1698431365
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1698431365
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1698431365
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1698431365
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1698431365
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1698431365
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1698431365
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1698431365
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1698431365
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1698431365
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1698431365
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1698431365
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1698431365
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1698431365
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1698431365
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1698431365
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1698431365
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1698431365
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1698431365
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1698431365
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1698431365
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1698431365
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1698431365
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1698431365
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1698431365
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1698431365
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1698431365
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1698431365
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1698431365
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1698431365
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1698431365
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1698431365
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1698431365
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1698431365
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1698431365
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1698431365
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1698431365
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1698431365
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1698431365
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1698431365
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1698431365
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1698431365
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1698431365
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1698431365
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1698431365
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1698431365
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1698431365
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1698431365
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1698431365
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1698431365
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1698431365
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1698431365
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1698431365
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1698431365
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1698431365
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1698431365
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1698431365
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1698431365
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1698431365
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1698431365
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1698431365
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1698431365
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1698431365
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1698431365
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1698431365
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1698431365
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1698431365
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1698431365
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1698431365
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1698431365
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1698431365
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1698431365
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1698431365
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1698431365
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1698431365
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1698431365
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1698431365
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1698431365
transform 1 0 24288 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 CLK_EXT
port 0 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 CLK_PLL
port 1 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 CLK_SR
port 2 nsew signal input
flabel metal3 s 27188 18504 27988 18624 0 FreeSans 480 0 0 0 Data_SR
port 3 nsew signal input
flabel metal2 s 24398 29332 24454 30132 0 FreeSans 224 90 0 0 NMOS1_PS1
port 4 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 NMOS1_PS2
port 5 nsew signal tristate
flabel metal2 s 10414 29332 10470 30132 0 FreeSans 224 90 0 0 NMOS2_PS1
port 6 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 NMOS2_PS2
port 7 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 NMOS_PS3
port 8 nsew signal tristate
flabel metal2 s 3422 29332 3478 30132 0 FreeSans 224 90 0 0 PMOS1_PS1
port 9 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 PMOS1_PS2
port 10 nsew signal tristate
flabel metal2 s 17406 29332 17462 30132 0 FreeSans 224 90 0 0 PMOS2_PS1
port 11 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 PMOS2_PS2
port 12 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 PMOS_PS3
port 13 nsew signal tristate
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 RST
port 14 nsew signal input
flabel metal3 s 27188 25848 27988 25968 0 FreeSans 480 0 0 0 SIGNAL_OUTPUT
port 15 nsew signal tristate
flabel metal4 s 4823 2128 5143 27792 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 11262 2128 11582 27792 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 17701 2128 18021 27792 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 24140 2128 24460 27792 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 5872 26912 6192 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 12264 26912 12584 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 18656 26912 18976 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 25048 26912 25368 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 4163 2128 4483 27792 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 10602 2128 10922 27792 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 17041 2128 17361 27792 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 23480 2128 23800 27792 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 5212 26912 5532 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 11604 26912 11924 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 17996 26912 18316 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 24388 26912 24708 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 d1[0]
port 18 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 d1[1]
port 19 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 d1[2]
port 20 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 d1[3]
port 21 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 d1[4]
port 22 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 d1[5]
port 23 nsew signal input
flabel metal3 s 27188 11160 27988 11280 0 FreeSans 480 0 0 0 d2[0]
port 24 nsew signal input
flabel metal3 s 27188 3816 27988 3936 0 FreeSans 480 0 0 0 d2[1]
port 25 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 d2[2]
port 26 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 d2[3]
port 27 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 d2[4]
port 28 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 d2[5]
port 29 nsew signal input
rlabel metal1 13984 27200 13984 27200 0 VGND
rlabel metal1 13984 27744 13984 27744 0 VPWR
rlabel metal2 2300 20740 2300 20740 0 CLK_EXT
rlabel metal1 2116 12206 2116 12206 0 CLK_PLL
rlabel metal1 10810 16524 10810 16524 0 CLK_SR
rlabel metal2 26542 18649 26542 18649 0 Data_SR
rlabel metal2 13110 13923 13110 13923 0 Dead_Time_Generator_inst_1.clk
rlabel metal1 7912 12818 7912 12818 0 Dead_Time_Generator_inst_1.count_dt\[0\]
rlabel metal1 7176 13498 7176 13498 0 Dead_Time_Generator_inst_1.count_dt\[1\]
rlabel metal1 7452 15334 7452 15334 0 Dead_Time_Generator_inst_1.count_dt\[2\]
rlabel metal2 7314 16286 7314 16286 0 Dead_Time_Generator_inst_1.count_dt\[3\]
rlabel metal2 9430 13634 9430 13634 0 Dead_Time_Generator_inst_1.count_dt\[4\]
rlabel via2 15134 12733 15134 12733 0 Dead_Time_Generator_inst_1.dt\[0\]
rlabel metal1 22494 13872 22494 13872 0 Dead_Time_Generator_inst_1.dt\[1\]
rlabel metal1 23092 13362 23092 13362 0 Dead_Time_Generator_inst_1.dt\[2\]
rlabel metal1 14122 13362 14122 13362 0 Dead_Time_Generator_inst_1.dt\[3\]
rlabel metal1 16422 13226 16422 13226 0 Dead_Time_Generator_inst_1.dt\[4\]
rlabel metal2 9890 16388 9890 16388 0 Dead_Time_Generator_inst_1.go
rlabel metal1 3220 16490 3220 16490 0 Dead_Time_Generator_inst_2.count_dt\[0\]
rlabel metal1 3726 14450 3726 14450 0 Dead_Time_Generator_inst_2.count_dt\[1\]
rlabel metal1 5106 16082 5106 16082 0 Dead_Time_Generator_inst_2.count_dt\[2\]
rlabel metal2 3266 13940 3266 13940 0 Dead_Time_Generator_inst_2.count_dt\[3\]
rlabel metal1 3818 13838 3818 13838 0 Dead_Time_Generator_inst_2.count_dt\[4\]
rlabel metal1 7636 17306 7636 17306 0 Dead_Time_Generator_inst_2.go
rlabel metal1 23598 14824 23598 14824 0 Dead_Time_Generator_inst_3.count_dt\[0\]
rlabel metal2 22862 15164 22862 15164 0 Dead_Time_Generator_inst_3.count_dt\[1\]
rlabel metal2 25070 14008 25070 14008 0 Dead_Time_Generator_inst_3.count_dt\[2\]
rlabel metal1 25254 13940 25254 13940 0 Dead_Time_Generator_inst_3.count_dt\[3\]
rlabel metal1 24794 12784 24794 12784 0 Dead_Time_Generator_inst_3.count_dt\[4\]
rlabel metal1 13478 17578 13478 17578 0 Dead_Time_Generator_inst_3.go
rlabel metal1 22034 10132 22034 10132 0 Dead_Time_Generator_inst_4.count_dt\[0\]
rlabel metal1 23184 9486 23184 9486 0 Dead_Time_Generator_inst_4.count_dt\[1\]
rlabel metal1 23644 9350 23644 9350 0 Dead_Time_Generator_inst_4.count_dt\[2\]
rlabel metal2 22770 9044 22770 9044 0 Dead_Time_Generator_inst_4.count_dt\[3\]
rlabel metal1 25668 11118 25668 11118 0 Dead_Time_Generator_inst_4.count_dt\[4\]
rlabel metal1 13018 16558 13018 16558 0 Dead_Time_Generator_inst_4.go
rlabel via1 24886 27557 24886 27557 0 NMOS1_PS1
rlabel metal2 17894 1095 17894 1095 0 NMOS1_PS2
rlabel metal1 10534 27574 10534 27574 0 NMOS2_PS1
rlabel metal2 9982 1554 9982 1554 0 NMOS2_PS2
rlabel metal2 25806 1520 25806 1520 0 NMOS_PS3
rlabel metal1 3680 27574 3680 27574 0 PMOS1_PS1
rlabel metal2 6026 1554 6026 1554 0 PMOS1_PS2
rlabel metal1 17618 27574 17618 27574 0 PMOS2_PS1
rlabel metal2 13938 1554 13938 1554 0 PMOS2_PS2
rlabel metal2 21850 1520 21850 1520 0 PMOS_PS3
rlabel metal3 820 23732 820 23732 0 RST
rlabel metal2 26174 26163 26174 26163 0 SIGNAL_OUTPUT
rlabel metal2 19550 19108 19550 19108 0 Shift_Register_Inst.data_out\[10\]
rlabel metal1 20194 18394 20194 18394 0 Shift_Register_Inst.data_out\[11\]
rlabel metal1 17480 20366 17480 20366 0 Shift_Register_Inst.data_out\[12\]
rlabel metal1 11592 16082 11592 16082 0 Shift_Register_Inst.data_out\[13\]
rlabel metal1 10810 12750 10810 12750 0 Shift_Register_Inst.data_out\[14\]
rlabel metal1 13570 17238 13570 17238 0 Shift_Register_Inst.data_out\[15\]
rlabel metal2 12834 13872 12834 13872 0 Shift_Register_Inst.data_out\[16\]
rlabel metal1 14168 14382 14168 14382 0 Shift_Register_Inst.data_out\[17\]
rlabel metal1 12788 22610 12788 22610 0 Shift_Register_Inst.data_out\[5\]
rlabel metal1 13110 22576 13110 22576 0 Shift_Register_Inst.data_out\[6\]
rlabel metal2 14214 10506 14214 10506 0 Shift_Register_Inst.data_out\[7\]
rlabel metal1 13616 10030 13616 10030 0 Shift_Register_Inst.data_out\[8\]
rlabel metal1 18538 18734 18538 18734 0 Shift_Register_Inst.data_out\[9\]
rlabel metal2 20654 13056 20654 13056 0 Shift_Register_Inst.shift_state\[0\]
rlabel metal2 21022 15266 21022 15266 0 Shift_Register_Inst.shift_state\[1\]
rlabel metal1 19550 16660 19550 16660 0 Shift_Register_Inst.shift_state\[2\]
rlabel metal1 17388 14382 17388 14382 0 Shift_Register_Inst.shift_state\[3\]
rlabel metal1 21206 16014 21206 16014 0 Shift_Register_Inst.shift_state\[4\]
rlabel metal1 20700 21998 20700 21998 0 Signal_Generator_1_0phase_inst.count\[0\]
rlabel metal1 22218 22984 22218 22984 0 Signal_Generator_1_0phase_inst.count\[1\]
rlabel metal1 17112 21522 17112 21522 0 Signal_Generator_1_0phase_inst.count\[2\]
rlabel metal2 18722 21930 18722 21930 0 Signal_Generator_1_0phase_inst.count\[3\]
rlabel metal1 19182 23494 19182 23494 0 Signal_Generator_1_0phase_inst.count\[4\]
rlabel metal2 18262 23919 18262 23919 0 Signal_Generator_1_0phase_inst.count\[5\]
rlabel metal2 23322 24412 23322 24412 0 Signal_Generator_1_0phase_inst.direction
rlabel metal2 7682 24582 7682 24582 0 Signal_Generator_1_180phase_inst.count\[0\]
rlabel metal1 7544 25806 7544 25806 0 Signal_Generator_1_180phase_inst.count\[1\]
rlabel metal2 8142 23970 8142 23970 0 Signal_Generator_1_180phase_inst.count\[2\]
rlabel metal2 8234 23698 8234 23698 0 Signal_Generator_1_180phase_inst.count\[3\]
rlabel via2 9338 23749 9338 23749 0 Signal_Generator_1_180phase_inst.count\[4\]
rlabel metal1 3818 24174 3818 24174 0 Signal_Generator_1_180phase_inst.count\[5\]
rlabel metal1 5106 25262 5106 25262 0 Signal_Generator_1_180phase_inst.direction
rlabel metal2 8234 21114 8234 21114 0 Signal_Generator_1_270phase_inst.count\[0\]
rlabel metal2 5198 18564 5198 18564 0 Signal_Generator_1_270phase_inst.count\[1\]
rlabel metal2 6854 20621 6854 20621 0 Signal_Generator_1_270phase_inst.count\[2\]
rlabel metal1 8426 21862 8426 21862 0 Signal_Generator_1_270phase_inst.count\[3\]
rlabel metal1 3496 20502 3496 20502 0 Signal_Generator_1_270phase_inst.count\[4\]
rlabel metal1 5060 21318 5060 21318 0 Signal_Generator_1_270phase_inst.count\[5\]
rlabel metal1 3312 19346 3312 19346 0 Signal_Generator_1_270phase_inst.direction
rlabel metal2 15226 23188 15226 23188 0 Signal_Generator_1_90phase_inst.count\[0\]
rlabel metal1 15226 26554 15226 26554 0 Signal_Generator_1_90phase_inst.count\[1\]
rlabel metal1 13432 24582 13432 24582 0 Signal_Generator_1_90phase_inst.count\[2\]
rlabel metal1 13938 24888 13938 24888 0 Signal_Generator_1_90phase_inst.count\[3\]
rlabel metal2 12926 24582 12926 24582 0 Signal_Generator_1_90phase_inst.count\[4\]
rlabel metal1 12512 24582 12512 24582 0 Signal_Generator_1_90phase_inst.count\[5\]
rlabel metal1 17342 26928 17342 26928 0 Signal_Generator_1_90phase_inst.direction
rlabel metal1 6302 2414 6302 2414 0 Signal_Generator_2_0phase_inst.count\[0\]
rlabel metal1 5612 2822 5612 2822 0 Signal_Generator_2_0phase_inst.count\[1\]
rlabel metal2 7406 3196 7406 3196 0 Signal_Generator_2_0phase_inst.count\[2\]
rlabel metal2 7498 6154 7498 6154 0 Signal_Generator_2_0phase_inst.count\[3\]
rlabel metal1 5474 7344 5474 7344 0 Signal_Generator_2_0phase_inst.count\[4\]
rlabel metal1 5658 6732 5658 6732 0 Signal_Generator_2_0phase_inst.count\[5\]
rlabel metal2 4462 6783 4462 6783 0 Signal_Generator_2_0phase_inst.direction
rlabel via1 20102 7939 20102 7939 0 Signal_Generator_2_180phase_inst.count\[0\]
rlabel metal1 15962 7174 15962 7174 0 Signal_Generator_2_180phase_inst.count\[1\]
rlabel metal2 20194 7004 20194 7004 0 Signal_Generator_2_180phase_inst.count\[2\]
rlabel metal1 19964 7922 19964 7922 0 Signal_Generator_2_180phase_inst.count\[3\]
rlabel metal1 17526 8364 17526 8364 0 Signal_Generator_2_180phase_inst.count\[4\]
rlabel metal1 16123 9350 16123 9350 0 Signal_Generator_2_180phase_inst.count\[5\]
rlabel metal2 20838 5542 20838 5542 0 Signal_Generator_2_180phase_inst.direction
rlabel metal1 11776 10234 11776 10234 0 Signal_Generator_2_270phase_inst.count\[0\]
rlabel metal2 8602 9180 8602 9180 0 Signal_Generator_2_270phase_inst.count\[1\]
rlabel metal1 11408 10574 11408 10574 0 Signal_Generator_2_270phase_inst.count\[2\]
rlabel metal1 12956 8874 12956 8874 0 Signal_Generator_2_270phase_inst.count\[3\]
rlabel metal1 13386 8942 13386 8942 0 Signal_Generator_2_270phase_inst.count\[4\]
rlabel metal2 6210 9112 6210 9112 0 Signal_Generator_2_270phase_inst.count\[5\]
rlabel metal2 7774 9792 7774 9792 0 Signal_Generator_2_270phase_inst.direction
rlabel metal1 11132 4046 11132 4046 0 Signal_Generator_2_90phase_inst.count\[0\]
rlabel metal1 14122 5032 14122 5032 0 Signal_Generator_2_90phase_inst.count\[1\]
rlabel metal1 13524 5202 13524 5202 0 Signal_Generator_2_90phase_inst.count\[2\]
rlabel metal1 14053 5814 14053 5814 0 Signal_Generator_2_90phase_inst.count\[3\]
rlabel metal1 14904 3910 14904 3910 0 Signal_Generator_2_90phase_inst.count\[4\]
rlabel metal1 15364 4182 15364 4182 0 Signal_Generator_2_90phase_inst.count\[5\]
rlabel metal1 16974 4692 16974 4692 0 Signal_Generator_2_90phase_inst.direction
rlabel metal1 16698 22066 16698 22066 0 _0000_
rlabel metal2 22310 23324 22310 23324 0 _0001_
rlabel metal2 22126 22814 22126 22814 0 _0002_
rlabel metal1 20056 22542 20056 22542 0 _0003_
rlabel metal2 19458 25534 19458 25534 0 _0004_
rlabel metal1 19780 25466 19780 25466 0 _0005_
rlabel metal2 22218 24276 22218 24276 0 _0006_
rlabel metal2 10258 24480 10258 24480 0 _0007_
rlabel metal1 4278 26350 4278 26350 0 _0008_
rlabel metal2 7314 26554 7314 26554 0 _0009_
rlabel metal2 6762 24140 6762 24140 0 _0010_
rlabel metal2 3726 24412 3726 24412 0 _0011_
rlabel metal1 1978 24718 1978 24718 0 _0012_
rlabel metal1 3680 26214 3680 26214 0 _0013_
rlabel metal1 6854 20026 6854 20026 0 _0014_
rlabel metal1 2691 18326 2691 18326 0 _0015_
rlabel metal1 6164 19278 6164 19278 0 _0016_
rlabel metal1 5888 21658 5888 21658 0 _0017_
rlabel metal1 2231 21454 2231 21454 0 _0018_
rlabel metal2 2990 21420 2990 21420 0 _0019_
rlabel metal1 3450 19278 3450 19278 0 _0020_
rlabel metal1 13754 23086 13754 23086 0 _0021_
rlabel metal1 16882 25670 16882 25670 0 _0022_
rlabel metal2 16882 24106 16882 24106 0 _0023_
rlabel metal1 13662 25806 13662 25806 0 _0024_
rlabel metal1 11362 25670 11362 25670 0 _0025_
rlabel metal1 11500 26010 11500 26010 0 _0026_
rlabel metal1 16606 25874 16606 25874 0 _0027_
rlabel metal2 8510 3604 8510 3604 0 _0028_
rlabel metal2 4002 3434 4002 3434 0 _0029_
rlabel metal2 6946 3298 6946 3298 0 _0030_
rlabel metal1 6440 4658 6440 4658 0 _0031_
rlabel metal1 3726 6834 3726 6834 0 _0032_
rlabel metal1 3864 6222 3864 6222 0 _0033_
rlabel metal2 4278 4352 4278 4352 0 _0034_
rlabel metal2 16330 6596 16330 6596 0 _0035_
rlabel metal1 19228 4114 19228 4114 0 _0036_
rlabel metal2 21022 7004 21022 7004 0 _0037_
rlabel metal2 19826 8228 19826 8228 0 _0038_
rlabel metal1 17848 9146 17848 9146 0 _0039_
rlabel metal1 16100 8602 16100 8602 0 _0040_
rlabel via1 19366 5219 19366 5219 0 _0041_
rlabel metal2 9982 10472 9982 10472 0 _0042_
rlabel metal2 5382 10778 5382 10778 0 _0043_
rlabel metal1 8556 10234 8556 10234 0 _0044_
rlabel metal1 10074 9350 10074 9350 0 _0045_
rlabel metal1 1886 9928 1886 9928 0 _0046_
rlabel metal1 3496 9486 3496 9486 0 _0047_
rlabel metal1 4554 10710 4554 10710 0 _0048_
rlabel metal1 9706 2958 9706 2958 0 _0049_
rlabel metal2 10442 3740 10442 3740 0 _0050_
rlabel metal1 14674 3570 14674 3570 0 _0051_
rlabel metal1 15134 4794 15134 4794 0 _0052_
rlabel metal2 17710 3706 17710 3706 0 _0053_
rlabel metal2 16974 3774 16974 3774 0 _0054_
rlabel metal2 10534 4828 10534 4828 0 _0055_
rlabel metal2 13570 13736 13570 13736 0 _0056_
rlabel metal1 12979 13226 12979 13226 0 _0057_
rlabel metal2 13110 15912 13110 15912 0 _0058_
rlabel metal1 11224 12954 11224 12954 0 _0059_
rlabel metal2 11270 15640 11270 15640 0 _0060_
rlabel metal1 18676 20026 18676 20026 0 _0061_
rlabel metal2 20010 19992 20010 19992 0 _0062_
rlabel metal2 20470 19176 20470 19176 0 _0063_
rlabel metal2 18906 19176 18906 19176 0 _0064_
rlabel metal1 13156 10778 13156 10778 0 _0065_
rlabel metal2 14582 10676 14582 10676 0 _0066_
rlabel metal1 15272 21658 15272 21658 0 _0067_
rlabel metal1 13708 21046 13708 21046 0 _0068_
rlabel metal2 16790 12002 16790 12002 0 _0069_
rlabel metal1 18860 12070 18860 12070 0 _0070_
rlabel metal2 20102 12002 20102 12002 0 _0071_
rlabel metal2 19642 10914 19642 10914 0 _0072_
rlabel metal1 19964 12954 19964 12954 0 _0073_
rlabel metal2 20930 15198 20930 15198 0 _0074_
rlabel metal1 20523 17238 20523 17238 0 _0075_
rlabel metal1 16744 16966 16744 16966 0 _0076_
rlabel metal2 20378 16286 20378 16286 0 _0077_
rlabel metal1 22448 24378 22448 24378 0 _0078_
rlabel metal1 17618 22066 17618 22066 0 _0079_
rlabel metal1 22724 23494 22724 23494 0 _0080_
rlabel metal2 22678 22372 22678 22372 0 _0081_
rlabel metal1 19925 22678 19925 22678 0 _0082_
rlabel metal2 19642 26146 19642 26146 0 _0083_
rlabel metal2 18998 26792 18998 26792 0 _0084_
rlabel metal2 18078 26078 18078 26078 0 _0085_
rlabel metal1 14444 23494 14444 23494 0 _0086_
rlabel metal2 16882 26520 16882 26520 0 _0087_
rlabel metal2 16330 23256 16330 23256 0 _0088_
rlabel metal2 14766 26078 14766 26078 0 _0089_
rlabel metal2 10350 26520 10350 26520 0 _0090_
rlabel metal2 12098 26520 12098 26520 0 _0091_
rlabel metal1 4515 25942 4515 25942 0 _0092_
rlabel metal1 9844 25466 9844 25466 0 _0093_
rlabel metal1 5152 26010 5152 26010 0 _0094_
rlabel metal1 8326 26323 8326 26323 0 _0095_
rlabel metal2 7130 23528 7130 23528 0 _0096_
rlabel metal2 2806 23970 2806 23970 0 _0097_
rlabel metal1 3312 24378 3312 24378 0 _0098_
rlabel metal1 2645 19414 2645 19414 0 _0099_
rlabel metal2 7314 20264 7314 20264 0 _0100_
rlabel metal2 3910 18462 3910 18462 0 _0101_
rlabel metal2 6946 19176 6946 19176 0 _0102_
rlabel metal1 7176 21658 7176 21658 0 _0103_
rlabel metal2 2806 21692 2806 21692 0 _0104_
rlabel metal2 2530 21352 2530 21352 0 _0105_
rlabel metal1 4002 3366 4002 3366 0 _0106_
rlabel metal2 8878 3672 8878 3672 0 _0107_
rlabel metal1 4784 3978 4784 3978 0 _0108_
rlabel metal1 8004 3162 8004 3162 0 _0109_
rlabel metal1 8103 4522 8103 4522 0 _0110_
rlabel metal1 2997 6698 2997 6698 0 _0111_
rlabel metal1 3687 6358 3687 6358 0 _0112_
rlabel metal1 9660 3706 9660 3706 0 _0113_
rlabel metal1 9706 2618 9706 2618 0 _0114_
rlabel metal1 11553 3434 11553 3434 0 _0115_
rlabel metal2 14858 3298 14858 3298 0 _0116_
rlabel metal2 15042 5848 15042 5848 0 _0117_
rlabel metal1 17395 3434 17395 3434 0 _0118_
rlabel metal2 18538 3230 18538 3230 0 _0119_
rlabel metal2 20010 4760 20010 4760 0 _0120_
rlabel metal2 16974 6562 16974 6562 0 _0121_
rlabel metal1 20523 4182 20523 4182 0 _0122_
rlabel metal2 21942 6562 21942 6562 0 _0123_
rlabel metal2 20562 8670 20562 8670 0 _0124_
rlabel metal2 16698 9384 16698 9384 0 _0125_
rlabel metal1 15640 9146 15640 9146 0 _0126_
rlabel metal1 3273 10710 3273 10710 0 _0127_
rlabel metal1 11231 9962 11231 9962 0 _0128_
rlabel metal2 6486 10914 6486 10914 0 _0129_
rlabel metal1 10350 9622 10350 9622 0 _0130_
rlabel metal2 12466 9792 12466 9792 0 _0131_
rlabel metal1 2852 9146 2852 9146 0 _0132_
rlabel metal2 3726 10030 3726 10030 0 _0133_
rlabel metal1 16054 11322 16054 11322 0 _0134_
rlabel metal2 12190 13396 12190 13396 0 _0135_
rlabel metal1 11040 13226 11040 13226 0 _0136_
rlabel metal2 12374 15844 12374 15844 0 _0137_
rlabel metal2 11086 13294 11086 13294 0 _0138_
rlabel metal2 10534 15640 10534 15640 0 _0139_
rlabel metal2 18446 20196 18446 20196 0 _0140_
rlabel metal1 19550 19720 19550 19720 0 _0141_
rlabel metal2 20102 19108 20102 19108 0 _0142_
rlabel metal1 17848 19278 17848 19278 0 _0143_
rlabel metal2 12374 11356 12374 11356 0 _0144_
rlabel metal1 14858 10778 14858 10778 0 _0145_
rlabel metal2 15686 21794 15686 21794 0 _0146_
rlabel metal1 13570 21114 13570 21114 0 _0147_
rlabel metal1 15870 12682 15870 12682 0 _0148_
rlabel metal1 17710 11798 17710 11798 0 _0149_
rlabel metal1 19136 11322 19136 11322 0 _0150_
rlabel metal1 19458 11186 19458 11186 0 _0151_
rlabel metal1 19366 13226 19366 13226 0 _0152_
rlabel metal1 19458 14586 19458 14586 0 _0153_
rlabel metal2 19090 17306 19090 17306 0 _0154_
rlabel metal2 15042 15844 15042 15844 0 _0155_
rlabel metal1 19320 15674 19320 15674 0 _0156_
rlabel metal1 21298 12206 21298 12206 0 _0157_
rlabel via1 10078 13294 10078 13294 0 _0158_
rlabel metal1 6297 13294 6297 13294 0 _0159_
rlabel metal1 5561 15402 5561 15402 0 _0160_
rlabel via1 6573 16490 6573 16490 0 _0161_
rlabel metal1 7447 17170 7447 17170 0 _0162_
rlabel metal1 16054 12614 16054 12614 0 _0163_
rlabel metal1 2300 15674 2300 15674 0 _0164_
rlabel metal1 1778 16150 1778 16150 0 _0165_
rlabel via1 4089 16558 4089 16558 0 _0166_
rlabel metal1 1962 13226 1962 13226 0 _0167_
rlabel metal2 3358 13532 3358 13532 0 _0168_
rlabel metal2 8602 15878 8602 15878 0 _0169_
rlabel metal2 21666 16082 21666 16082 0 _0170_
rlabel metal1 23240 15470 23240 15470 0 _0171_
rlabel metal1 24973 15470 24973 15470 0 _0172_
rlabel metal1 24548 14314 24548 14314 0 _0173_
rlabel metal1 24932 12954 24932 12954 0 _0174_
rlabel metal1 5198 16762 5198 16762 0 _0175_
rlabel metal2 21298 9826 21298 9826 0 _0176_
rlabel metal2 22494 8738 22494 8738 0 _0177_
rlabel metal1 25571 9962 25571 9962 0 _0178_
rlabel viali 23878 8534 23878 8534 0 _0179_
rlabel metal1 24502 10710 24502 10710 0 _0180_
rlabel metal2 21666 17102 21666 17102 0 _0181_
rlabel metal2 14490 21182 14490 21182 0 _0182_
rlabel metal1 17434 13872 17434 13872 0 _0183_
rlabel metal2 15042 12954 15042 12954 0 _0184_
rlabel metal1 15640 12818 15640 12818 0 _0185_
rlabel metal1 16422 16762 16422 16762 0 _0186_
rlabel metal2 16882 14688 16882 14688 0 _0187_
rlabel metal1 18400 15130 18400 15130 0 _0188_
rlabel metal1 17342 16048 17342 16048 0 _0189_
rlabel metal1 14858 15470 14858 15470 0 _0190_
rlabel metal1 15134 15504 15134 15504 0 _0191_
rlabel metal1 17710 16082 17710 16082 0 _0192_
rlabel metal1 18078 16014 18078 16014 0 _0193_
rlabel metal1 18952 14586 18952 14586 0 _0194_
rlabel metal2 18630 13634 18630 13634 0 _0195_
rlabel metal1 18492 14042 18492 14042 0 _0196_
rlabel metal1 19228 14382 19228 14382 0 _0197_
rlabel metal1 18032 12750 18032 12750 0 _0198_
rlabel metal1 18308 11118 18308 11118 0 _0199_
rlabel metal2 19458 15504 19458 15504 0 _0200_
rlabel metal1 19136 12750 19136 12750 0 _0201_
rlabel metal2 18538 11866 18538 11866 0 _0202_
rlabel metal1 17894 14858 17894 14858 0 _0203_
rlabel metal2 17342 11900 17342 11900 0 _0204_
rlabel metal2 17986 14739 17986 14739 0 _0205_
rlabel metal1 15962 13362 15962 13362 0 _0206_
rlabel metal2 16146 12988 16146 12988 0 _0207_
rlabel metal2 9384 21862 9384 21862 0 _0208_
rlabel metal1 16376 16694 16376 16694 0 _0209_
rlabel metal1 12926 20876 12926 20876 0 _0210_
rlabel metal1 13984 22406 13984 22406 0 _0211_
rlabel via2 15410 17323 15410 17323 0 _0212_
rlabel metal1 15502 21488 15502 21488 0 _0213_
rlabel metal1 14444 10166 14444 10166 0 _0214_
rlabel metal1 14030 10642 14030 10642 0 _0215_
rlabel metal2 13754 10914 13754 10914 0 _0216_
rlabel metal1 16744 14246 16744 14246 0 _0217_
rlabel metal1 13432 11730 13432 11730 0 _0218_
rlabel metal2 18078 17612 18078 17612 0 _0219_
rlabel metal1 18078 18938 18078 18938 0 _0220_
rlabel metal2 19826 17612 19826 17612 0 _0221_
rlabel metal1 20148 18734 20148 18734 0 _0222_
rlabel metal1 19044 17306 19044 17306 0 _0223_
rlabel metal2 18998 19108 18998 19108 0 _0224_
rlabel metal2 16698 15266 16698 15266 0 _0225_
rlabel metal2 17526 17782 17526 17782 0 _0226_
rlabel metal1 18262 19856 18262 19856 0 _0227_
rlabel metal1 10304 19346 10304 19346 0 _0228_
rlabel metal2 15226 16184 15226 16184 0 _0229_
rlabel metal1 11086 16150 11086 16150 0 _0230_
rlabel metal2 13294 12818 13294 12818 0 _0231_
rlabel metal1 11638 12954 11638 12954 0 _0232_
rlabel metal1 14720 16014 14720 16014 0 _0233_
rlabel metal1 12834 15504 12834 15504 0 _0234_
rlabel metal2 14582 14246 14582 14246 0 _0235_
rlabel metal2 11730 14076 11730 14076 0 _0236_
rlabel metal1 15167 14042 15167 14042 0 _0237_
rlabel metal1 14398 13804 14398 13804 0 _0238_
rlabel metal1 12972 12818 12972 12818 0 _0239_
rlabel metal2 18538 22644 18538 22644 0 _0240_
rlabel metal1 19872 24174 19872 24174 0 _0241_
rlabel metal1 19136 24378 19136 24378 0 _0242_
rlabel metal1 20525 23018 20525 23018 0 _0243_
rlabel via1 19918 24854 19918 24854 0 _0244_
rlabel metal1 19504 23562 19504 23562 0 _0245_
rlabel metal1 21114 22406 21114 22406 0 _0246_
rlabel metal1 22586 23732 22586 23732 0 _0247_
rlabel metal1 22310 23630 22310 23630 0 _0248_
rlabel metal1 21344 22202 21344 22202 0 _0249_
rlabel metal1 21528 22542 21528 22542 0 _0250_
rlabel metal2 22126 23392 22126 23392 0 _0251_
rlabel metal1 18308 21658 18308 21658 0 _0252_
rlabel metal2 19734 23188 19734 23188 0 _0253_
rlabel metal2 19826 24276 19826 24276 0 _0254_
rlabel metal1 19182 22202 19182 22202 0 _0255_
rlabel metal1 19044 23018 19044 23018 0 _0256_
rlabel metal1 19182 24752 19182 24752 0 _0257_
rlabel metal1 19320 24786 19320 24786 0 _0258_
rlabel metal2 18814 24956 18814 24956 0 _0259_
rlabel metal1 19044 24650 19044 24650 0 _0260_
rlabel metal1 13064 25398 13064 25398 0 _0261_
rlabel metal2 12742 26010 12742 26010 0 _0262_
rlabel metal2 15778 25500 15778 25500 0 _0263_
rlabel metal1 13064 23698 13064 23698 0 _0264_
rlabel metal1 13792 24854 13792 24854 0 _0265_
rlabel metal1 13202 26928 13202 26928 0 _0266_
rlabel metal2 15962 25364 15962 25364 0 _0267_
rlabel metal1 15502 25262 15502 25262 0 _0268_
rlabel metal2 16054 25670 16054 25670 0 _0269_
rlabel metal1 16100 25942 16100 25942 0 _0270_
rlabel metal1 16606 25296 16606 25296 0 _0271_
rlabel metal1 15594 24752 15594 24752 0 _0272_
rlabel metal1 16284 24922 16284 24922 0 _0273_
rlabel metal1 12926 25874 12926 25874 0 _0274_
rlabel metal1 12696 25738 12696 25738 0 _0275_
rlabel metal2 13110 25772 13110 25772 0 _0276_
rlabel metal1 13018 24752 13018 24752 0 _0277_
rlabel metal2 13478 25602 13478 25602 0 _0278_
rlabel metal1 12190 24922 12190 24922 0 _0279_
rlabel metal1 11868 24922 11868 24922 0 _0280_
rlabel metal1 11592 25398 11592 25398 0 _0281_
rlabel metal2 11546 25602 11546 25602 0 _0282_
rlabel metal1 6026 24718 6026 24718 0 _0283_
rlabel metal1 5106 24786 5106 24786 0 _0284_
rlabel metal1 6670 24820 6670 24820 0 _0285_
rlabel metal1 6578 26350 6578 26350 0 _0286_
rlabel via1 4638 25126 4638 25126 0 _0287_
rlabel metal1 5980 24174 5980 24174 0 _0288_
rlabel metal1 7130 25772 7130 25772 0 _0289_
rlabel metal1 4186 26996 4186 26996 0 _0290_
rlabel metal2 3634 26554 3634 26554 0 _0291_
rlabel metal1 6808 25670 6808 25670 0 _0292_
rlabel metal1 7038 26554 7038 26554 0 _0293_
rlabel metal1 7176 27030 7176 27030 0 _0294_
rlabel metal2 6210 24548 6210 24548 0 _0295_
rlabel metal1 6762 24752 6762 24752 0 _0296_
rlabel metal1 6762 24038 6762 24038 0 _0297_
rlabel metal1 6762 24208 6762 24208 0 _0298_
rlabel metal1 6440 24378 6440 24378 0 _0299_
rlabel metal1 7590 24106 7590 24106 0 _0300_
rlabel metal1 4232 24378 4232 24378 0 _0301_
rlabel metal1 4094 23834 4094 23834 0 _0302_
rlabel metal1 4324 24854 4324 24854 0 _0303_
rlabel metal1 5060 24038 5060 24038 0 _0304_
rlabel metal1 4232 21046 4232 21046 0 _0305_
rlabel metal1 4508 20910 4508 20910 0 _0306_
rlabel viali 3713 21522 3713 21522 0 _0307_
rlabel metal1 4830 19822 4830 19822 0 _0308_
rlabel metal1 4600 21981 4600 21981 0 _0309_
rlabel metal1 4002 19346 4002 19346 0 _0310_
rlabel metal1 4784 19278 4784 19278 0 _0311_
rlabel metal2 3542 19516 3542 19516 0 _0312_
rlabel metal1 2852 19346 2852 19346 0 _0313_
rlabel metal1 5244 19278 5244 19278 0 _0314_
rlabel metal1 5428 18938 5428 18938 0 _0315_
rlabel metal1 5428 19414 5428 19414 0 _0316_
rlabel metal2 5566 21284 5566 21284 0 _0317_
rlabel metal2 5382 21692 5382 21692 0 _0318_
rlabel metal1 4554 21556 4554 21556 0 _0319_
rlabel metal1 4738 20944 4738 20944 0 _0320_
rlabel metal2 5198 21313 5198 21313 0 _0321_
rlabel metal1 3910 21624 3910 21624 0 _0322_
rlabel metal1 4048 20570 4048 20570 0 _0323_
rlabel metal1 3496 20570 3496 20570 0 _0324_
rlabel metal1 3634 21998 3634 21998 0 _0325_
rlabel metal2 6118 6596 6118 6596 0 _0326_
rlabel metal2 5934 6970 5934 6970 0 _0327_
rlabel metal1 4554 4080 4554 4080 0 _0328_
rlabel metal1 6348 3910 6348 3910 0 _0329_
rlabel metal2 5658 7684 5658 7684 0 _0330_
rlabel metal1 5106 4590 5106 4590 0 _0331_
rlabel metal1 5658 2618 5658 2618 0 _0332_
rlabel metal2 4462 4318 4462 4318 0 _0333_
rlabel metal1 4462 3910 4462 3910 0 _0334_
rlabel metal1 7038 2992 7038 2992 0 _0335_
rlabel metal1 5750 2958 5750 2958 0 _0336_
rlabel metal1 6394 3094 6394 3094 0 _0337_
rlabel metal2 6302 6324 6302 6324 0 _0338_
rlabel metal2 6026 6460 6026 6460 0 _0339_
rlabel metal1 5244 6290 5244 6290 0 _0340_
rlabel metal1 5106 6256 5106 6256 0 _0341_
rlabel metal1 5704 6358 5704 6358 0 _0342_
rlabel metal1 4370 6664 4370 6664 0 _0343_
rlabel metal1 4554 6766 4554 6766 0 _0344_
rlabel metal2 4738 7004 4738 7004 0 _0345_
rlabel metal1 4508 6426 4508 6426 0 _0346_
rlabel metal1 17342 3978 17342 3978 0 _0347_
rlabel metal2 17250 4284 17250 4284 0 _0348_
rlabel metal1 17181 4182 17181 4182 0 _0349_
rlabel metal1 13156 4522 13156 4522 0 _0350_
rlabel metal1 14477 4250 14477 4250 0 _0351_
rlabel metal1 13478 4216 13478 4216 0 _0352_
rlabel metal1 12926 3570 12926 3570 0 _0353_
rlabel metal1 11730 4114 11730 4114 0 _0354_
rlabel metal1 11588 4250 11588 4250 0 _0355_
rlabel metal1 13570 3536 13570 3536 0 _0356_
rlabel metal1 13202 4080 13202 4080 0 _0357_
rlabel metal2 13386 3706 13386 3706 0 _0358_
rlabel via2 15134 5219 15134 5219 0 _0359_
rlabel metal1 14674 4590 14674 4590 0 _0360_
rlabel metal2 15686 4284 15686 4284 0 _0361_
rlabel metal1 15134 4590 15134 4590 0 _0362_
rlabel metal1 14306 4624 14306 4624 0 _0363_
rlabel metal2 17802 4063 17802 4063 0 _0364_
rlabel metal1 18032 4114 18032 4114 0 _0365_
rlabel metal2 17434 4420 17434 4420 0 _0366_
rlabel metal1 18124 4250 18124 4250 0 _0367_
rlabel metal1 18032 8398 18032 8398 0 _0368_
rlabel metal1 19044 8466 19044 8466 0 _0369_
rlabel metal1 18400 8602 18400 8602 0 _0370_
rlabel metal1 20516 6834 20516 6834 0 _0371_
rlabel metal1 19964 8942 19964 8942 0 _0372_
rlabel metal1 20838 7854 20838 7854 0 _0373_
rlabel metal1 19734 6256 19734 6256 0 _0374_
rlabel metal2 19642 5882 19642 5882 0 _0375_
rlabel metal1 19274 5270 19274 5270 0 _0376_
rlabel metal2 20930 6732 20930 6732 0 _0377_
rlabel metal2 20562 7395 20562 7395 0 _0378_
rlabel metal1 20608 7446 20608 7446 0 _0379_
rlabel metal1 18354 7514 18354 7514 0 _0380_
rlabel metal1 19642 7888 19642 7888 0 _0381_
rlabel metal1 18446 7956 18446 7956 0 _0382_
rlabel metal1 20700 7378 20700 7378 0 _0383_
rlabel metal1 20516 7514 20516 7514 0 _0384_
rlabel metal2 18170 8432 18170 8432 0 _0385_
rlabel metal1 17710 8976 17710 8976 0 _0386_
rlabel metal1 18170 9044 18170 9044 0 _0387_
rlabel metal1 17710 8398 17710 8398 0 _0388_
rlabel metal2 4140 9350 4140 9350 0 _0389_
rlabel metal2 5198 10234 5198 10234 0 _0390_
rlabel metal1 8050 9928 8050 9928 0 _0391_
rlabel metal2 7130 9316 7130 9316 0 _0392_
rlabel metal1 4462 9588 4462 9588 0 _0393_
rlabel metal2 6854 10370 6854 10370 0 _0394_
rlabel metal1 7406 10132 7406 10132 0 _0395_
rlabel metal2 5934 10336 5934 10336 0 _0396_
rlabel metal1 5382 10608 5382 10608 0 _0397_
rlabel metal1 8142 10064 8142 10064 0 _0398_
rlabel metal2 7406 10064 7406 10064 0 _0399_
rlabel metal1 7912 10030 7912 10030 0 _0400_
rlabel metal1 8602 9996 8602 9996 0 _0401_
rlabel metal1 8234 9554 8234 9554 0 _0402_
rlabel metal2 6026 9520 6026 9520 0 _0403_
rlabel metal1 7958 9486 7958 9486 0 _0404_
rlabel metal2 7866 9758 7866 9758 0 _0405_
rlabel metal1 4646 9690 4646 9690 0 _0406_
rlabel metal1 4186 10064 4186 10064 0 _0407_
rlabel metal1 4508 9078 4508 9078 0 _0408_
rlabel metal2 4738 10030 4738 10030 0 _0409_
rlabel metal1 3174 12274 3174 12274 0 _0410_
rlabel metal2 13754 19550 13754 19550 0 _0411_
rlabel metal1 13524 18802 13524 18802 0 _0412_
rlabel metal1 14214 17272 14214 17272 0 _0413_
rlabel metal2 13570 17204 13570 17204 0 _0414_
rlabel metal1 14766 17170 14766 17170 0 _0415_
rlabel metal1 13478 18156 13478 18156 0 _0416_
rlabel metal2 13570 18122 13570 18122 0 _0417_
rlabel metal1 14674 18156 14674 18156 0 _0418_
rlabel metal2 9430 17476 9430 17476 0 _0419_
rlabel metal1 11086 17170 11086 17170 0 _0420_
rlabel metal1 9844 16762 9844 16762 0 _0421_
rlabel metal1 10672 16966 10672 16966 0 _0422_
rlabel metal2 11638 16932 11638 16932 0 _0423_
rlabel metal1 13892 17646 13892 17646 0 _0424_
rlabel metal1 15318 17612 15318 17612 0 _0425_
rlabel metal1 14168 18394 14168 18394 0 _0426_
rlabel metal1 10028 17850 10028 17850 0 _0427_
rlabel metal2 10534 18122 10534 18122 0 _0428_
rlabel metal1 17526 20774 17526 20774 0 _0429_
rlabel metal1 15916 18734 15916 18734 0 _0430_
rlabel metal2 17066 19601 17066 19601 0 _0431_
rlabel metal1 15870 18632 15870 18632 0 _0432_
rlabel metal1 15456 19958 15456 19958 0 _0433_
rlabel metal1 17020 19482 17020 19482 0 _0434_
rlabel metal2 16146 20128 16146 20128 0 _0435_
rlabel metal2 16514 20196 16514 20196 0 _0436_
rlabel metal1 15594 18292 15594 18292 0 _0437_
rlabel metal1 15272 18394 15272 18394 0 _0438_
rlabel metal1 15042 18666 15042 18666 0 _0439_
rlabel metal1 15502 18938 15502 18938 0 _0440_
rlabel metal1 17158 18768 17158 18768 0 _0441_
rlabel metal2 16514 19108 16514 19108 0 _0442_
rlabel metal1 16547 18394 16547 18394 0 _0443_
rlabel metal1 16652 18122 16652 18122 0 _0444_
rlabel metal1 15778 19210 15778 19210 0 _0445_
rlabel metal1 14674 10642 14674 10642 0 _0446_
rlabel metal2 16054 11186 16054 11186 0 _0447_
rlabel metal2 18814 20162 18814 20162 0 _0448_
rlabel metal2 20838 16320 20838 16320 0 _0449_
rlabel metal1 22586 21964 22586 21964 0 _0450_
rlabel metal2 23230 11526 23230 11526 0 _0451_
rlabel metal1 22586 11118 22586 11118 0 _0452_
rlabel metal2 22034 11526 22034 11526 0 _0453_
rlabel metal1 22862 11764 22862 11764 0 _0454_
rlabel metal2 22954 11492 22954 11492 0 _0455_
rlabel metal2 22678 11900 22678 11900 0 _0456_
rlabel metal1 23552 11730 23552 11730 0 _0457_
rlabel metal1 23828 11322 23828 11322 0 _0458_
rlabel metal1 24058 11594 24058 11594 0 _0459_
rlabel metal1 24380 11730 24380 11730 0 _0460_
rlabel metal2 21482 11866 21482 11866 0 _0461_
rlabel metal2 2254 5848 2254 5848 0 _0462_
rlabel metal1 14763 7854 14763 7854 0 _0463_
rlabel metal2 14858 8024 14858 8024 0 _0464_
rlabel metal2 15134 8330 15134 8330 0 _0465_
rlabel metal1 11822 7480 11822 7480 0 _0466_
rlabel metal1 8188 7310 8188 7310 0 _0467_
rlabel metal2 7498 7650 7498 7650 0 _0468_
rlabel metal1 9200 6834 9200 6834 0 _0469_
rlabel metal1 2507 7922 2507 7922 0 _0470_
rlabel metal1 14996 8058 14996 8058 0 _0471_
rlabel metal2 15226 7225 15226 7225 0 _0472_
rlabel metal2 8418 7548 8418 7548 0 _0473_
rlabel metal2 8326 7174 8326 7174 0 _0474_
rlabel metal2 8786 7582 8786 7582 0 _0475_
rlabel metal1 8786 7378 8786 7378 0 _0476_
rlabel metal1 9384 6970 9384 6970 0 _0477_
rlabel metal1 9430 5610 9430 5610 0 _0478_
rlabel metal2 13386 8160 13386 8160 0 _0479_
rlabel metal1 13294 8364 13294 8364 0 _0480_
rlabel metal1 13110 8534 13110 8534 0 _0481_
rlabel metal2 12926 7106 12926 7106 0 _0482_
rlabel via2 8970 6307 8970 6307 0 _0483_
rlabel metal1 10304 6290 10304 6290 0 _0484_
rlabel metal1 9706 5576 9706 5576 0 _0485_
rlabel metal2 13662 7072 13662 7072 0 _0486_
rlabel metal1 13662 6868 13662 6868 0 _0487_
rlabel metal2 12834 9214 12834 9214 0 _0488_
rlabel metal1 11638 5610 11638 5610 0 _0489_
rlabel metal1 8702 6426 8702 6426 0 _0490_
rlabel metal1 9890 6120 9890 6120 0 _0491_
rlabel metal1 10166 5848 10166 5848 0 _0492_
rlabel metal1 9660 6358 9660 6358 0 _0493_
rlabel metal1 10166 6086 10166 6086 0 _0494_
rlabel metal1 11776 7378 11776 7378 0 _0495_
rlabel metal1 11270 7174 11270 7174 0 _0496_
rlabel metal1 10258 6630 10258 6630 0 _0497_
rlabel metal2 12006 7786 12006 7786 0 _0498_
rlabel metal1 12282 7956 12282 7956 0 _0499_
rlabel metal2 12098 8330 12098 8330 0 _0500_
rlabel metal2 12466 7242 12466 7242 0 _0501_
rlabel metal1 12788 6698 12788 6698 0 _0502_
rlabel metal1 11454 7820 11454 7820 0 _0503_
rlabel metal1 11776 7854 11776 7854 0 _0504_
rlabel metal1 11454 6800 11454 6800 0 _0505_
rlabel metal1 11546 6732 11546 6732 0 _0506_
rlabel viali 9890 6767 9890 6767 0 _0507_
rlabel metal2 10718 6596 10718 6596 0 _0508_
rlabel metal1 10626 6800 10626 6800 0 _0509_
rlabel metal2 10350 7123 10350 7123 0 _0510_
rlabel metal2 9798 6970 9798 6970 0 _0511_
rlabel metal2 20746 7310 20746 7310 0 _0512_
rlabel metal1 23874 16014 23874 16014 0 _0513_
rlabel metal1 21988 12410 21988 12410 0 _0514_
rlabel metal2 14858 26724 14858 26724 0 _0515_
rlabel metal2 2438 20672 2438 20672 0 _0516_
rlabel metal1 9246 2414 9246 2414 0 _0517_
rlabel metal2 15226 4658 15226 4658 0 _0518_
rlabel metal2 11822 20230 11822 20230 0 _0519_
rlabel metal1 12236 22406 12236 22406 0 _0520_
rlabel metal2 11086 23698 11086 23698 0 _0521_
rlabel metal1 11684 22066 11684 22066 0 _0522_
rlabel metal1 11224 22202 11224 22202 0 _0523_
rlabel metal1 11546 20536 11546 20536 0 _0524_
rlabel metal1 10994 19890 10994 19890 0 _0525_
rlabel metal1 11592 19754 11592 19754 0 _0526_
rlabel metal1 10304 20026 10304 20026 0 _0527_
rlabel metal1 10580 19686 10580 19686 0 _0528_
rlabel metal1 9430 19380 9430 19380 0 _0529_
rlabel metal1 10120 18938 10120 18938 0 _0530_
rlabel metal1 9016 22610 9016 22610 0 _0531_
rlabel metal1 10994 22712 10994 22712 0 _0532_
rlabel metal2 11822 22916 11822 22916 0 _0533_
rlabel metal1 10718 19244 10718 19244 0 _0534_
rlabel metal2 9062 19380 9062 19380 0 _0535_
rlabel metal1 10488 22610 10488 22610 0 _0536_
rlabel metal2 13018 22848 13018 22848 0 _0537_
rlabel metal2 10994 23052 10994 23052 0 _0538_
rlabel metal1 10396 19822 10396 19822 0 _0539_
rlabel metal1 11270 19278 11270 19278 0 _0540_
rlabel metal2 9430 19754 9430 19754 0 _0541_
rlabel metal1 10810 20434 10810 20434 0 _0542_
rlabel metal2 9890 22338 9890 22338 0 _0543_
rlabel metal1 9706 22440 9706 22440 0 _0544_
rlabel metal1 9522 21862 9522 21862 0 _0545_
rlabel metal2 9706 22559 9706 22559 0 _0546_
rlabel metal1 10166 20536 10166 20536 0 _0547_
rlabel metal2 10994 21148 10994 21148 0 _0548_
rlabel via1 9969 20434 9969 20434 0 _0549_
rlabel metal1 10166 20944 10166 20944 0 _0550_
rlabel metal1 10074 20298 10074 20298 0 _0551_
rlabel metal1 9936 20230 9936 20230 0 _0552_
rlabel metal1 9568 20570 9568 20570 0 _0553_
rlabel metal1 9062 20570 9062 20570 0 _0554_
rlabel metal2 8694 20298 8694 20298 0 _0555_
rlabel metal1 8786 19890 8786 19890 0 _0556_
rlabel metal1 10074 19788 10074 19788 0 _0557_
rlabel metal2 8786 19516 8786 19516 0 _0558_
rlabel metal2 9522 19550 9522 19550 0 _0559_
rlabel metal1 9798 19346 9798 19346 0 _0560_
rlabel metal1 8418 15504 8418 15504 0 _0561_
rlabel metal1 8188 13294 8188 13294 0 _0562_
rlabel metal1 8326 12954 8326 12954 0 _0563_
rlabel metal1 7774 13158 7774 13158 0 _0564_
rlabel metal2 7498 13770 7498 13770 0 _0565_
rlabel metal1 8602 14042 8602 14042 0 _0566_
rlabel metal2 7774 14858 7774 14858 0 _0567_
rlabel metal2 8280 12580 8280 12580 0 _0568_
rlabel metal1 8556 12342 8556 12342 0 _0569_
rlabel metal1 8648 12750 8648 12750 0 _0570_
rlabel metal1 8740 12682 8740 12682 0 _0571_
rlabel metal2 8694 13532 8694 13532 0 _0572_
rlabel metal1 8188 14382 8188 14382 0 _0573_
rlabel metal2 8234 14110 8234 14110 0 _0574_
rlabel metal2 9798 14076 9798 14076 0 _0575_
rlabel metal1 7360 15470 7360 15470 0 _0576_
rlabel metal2 6670 14076 6670 14076 0 _0577_
rlabel metal1 5704 15130 5704 15130 0 _0578_
rlabel metal1 7682 16218 7682 16218 0 _0579_
rlabel metal1 9016 16626 9016 16626 0 _0580_
rlabel metal1 8280 17170 8280 17170 0 _0581_
rlabel metal2 5290 13804 5290 13804 0 _0582_
rlabel metal2 4922 13549 4922 13549 0 _0583_
rlabel metal2 5566 13668 5566 13668 0 _0584_
rlabel metal1 5520 12818 5520 12818 0 _0585_
rlabel metal1 5106 12682 5106 12682 0 _0586_
rlabel metal1 4554 13328 4554 13328 0 _0587_
rlabel metal1 4646 13498 4646 13498 0 _0588_
rlabel metal2 4738 13260 4738 13260 0 _0589_
rlabel metal1 4692 12410 4692 12410 0 _0590_
rlabel metal1 4554 12716 4554 12716 0 _0591_
rlabel metal1 4508 12818 4508 12818 0 _0592_
rlabel metal1 3558 15062 3558 15062 0 _0593_
rlabel metal1 3266 15368 3266 15368 0 _0594_
rlabel metal1 2990 15674 2990 15674 0 _0595_
rlabel metal1 2576 15470 2576 15470 0 _0596_
rlabel metal1 3680 14790 3680 14790 0 _0597_
rlabel metal2 3634 15776 3634 15776 0 _0598_
rlabel metal1 1426 16048 1426 16048 0 _0599_
rlabel metal2 3910 16422 3910 16422 0 _0600_
rlabel metal2 4140 13498 4140 13498 0 _0601_
rlabel metal2 2806 13974 2806 13974 0 _0602_
rlabel metal1 1656 13294 1656 13294 0 _0603_
rlabel metal1 22678 13906 22678 13906 0 _0604_
rlabel metal2 22218 14076 22218 14076 0 _0605_
rlabel metal1 22724 13974 22724 13974 0 _0606_
rlabel metal1 23644 13906 23644 13906 0 _0607_
rlabel metal1 22816 14042 22816 14042 0 _0608_
rlabel metal1 23046 14382 23046 14382 0 _0609_
rlabel metal1 22770 13498 22770 13498 0 _0610_
rlabel metal1 23782 13328 23782 13328 0 _0611_
rlabel metal2 23874 13838 23874 13838 0 _0612_
rlabel metal1 23874 12954 23874 12954 0 _0613_
rlabel metal1 24518 12954 24518 12954 0 _0614_
rlabel metal1 23322 16694 23322 16694 0 _0615_
rlabel metal1 23644 16626 23644 16626 0 _0616_
rlabel metal1 22494 16966 22494 16966 0 _0617_
rlabel metal1 24150 15130 24150 15130 0 _0618_
rlabel metal2 24058 16252 24058 16252 0 _0619_
rlabel metal1 25116 15130 25116 15130 0 _0620_
rlabel metal2 24886 14314 24886 14314 0 _0621_
rlabel metal2 24242 14586 24242 14586 0 _0622_
rlabel metal2 23046 9724 23046 9724 0 _0623_
rlabel metal1 22264 10234 22264 10234 0 _0624_
rlabel metal1 21482 9588 21482 9588 0 _0625_
rlabel metal1 21390 8908 21390 8908 0 _0626_
rlabel metal2 22218 9248 22218 9248 0 _0627_
rlabel metal2 22678 8636 22678 8636 0 _0628_
rlabel metal2 25162 9622 25162 9622 0 _0629_
rlabel metal1 25500 9622 25500 9622 0 _0630_
rlabel metal2 25346 9860 25346 9860 0 _0631_
rlabel metal2 24058 10064 24058 10064 0 _0632_
rlabel metal1 23460 9146 23460 9146 0 _0633_
rlabel metal1 23414 9078 23414 9078 0 _0634_
rlabel metal1 16008 15470 16008 15470 0 clknet_0_CLK_SR
rlabel metal2 14398 16218 14398 16218 0 clknet_0_Dead_Time_Generator_inst_1.clk
rlabel metal1 19320 13362 19320 13362 0 clknet_1_0__leaf_CLK_SR
rlabel metal2 15962 21794 15962 21794 0 clknet_1_1__leaf_CLK_SR
rlabel metal2 4186 6494 4186 6494 0 clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 2300 13294 2300 13294 0 clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 19228 4658 19228 4658 0 clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 24656 13362 24656 13362 0 clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 1932 18258 1932 18258 0 clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 2024 24786 2024 24786 0 clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 23920 15538 23920 15538 0 clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 13386 24208 13386 24208 0 clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal3 1050 10676 1050 10676 0 d1[0]
rlabel metal3 1050 12852 1050 12852 0 d1[1]
rlabel metal3 1050 15028 1050 15028 0 d1[2]
rlabel metal3 820 17204 820 17204 0 d1[3]
rlabel metal3 820 19380 820 19380 0 d1[4]
rlabel metal3 820 21556 820 21556 0 d1[5]
rlabel metal2 26542 11475 26542 11475 0 d2[0]
rlabel metal2 26542 3995 26542 3995 0 d2[1]
rlabel metal3 820 1972 820 1972 0 d2[2]
rlabel metal3 820 4148 820 4148 0 d2[3]
rlabel metal3 820 6324 820 6324 0 d2[4]
rlabel metal3 820 8500 820 8500 0 d2[5]
rlabel metal2 19458 18462 19458 18462 0 net1
rlabel metal2 26358 4828 26358 4828 0 net10
rlabel metal1 2024 2618 2024 2618 0 net11
rlabel metal2 1610 4998 1610 4998 0 net12
rlabel metal1 1886 6290 1886 6290 0 net13
rlabel metal2 2162 8330 2162 8330 0 net14
rlabel metal2 24610 23970 24610 23970 0 net15
rlabel metal1 16974 2414 16974 2414 0 net16
rlabel metal2 14490 20094 14490 20094 0 net17
rlabel metal1 10810 2414 10810 2414 0 net18
rlabel metal1 25990 2448 25990 2448 0 net19
rlabel metal1 2254 23800 2254 23800 0 net2
rlabel metal2 15870 20077 15870 20077 0 net20
rlabel metal1 6762 2448 6762 2448 0 net21
rlabel metal1 16698 19448 16698 19448 0 net22
rlabel metal1 14398 2414 14398 2414 0 net23
rlabel metal2 15962 18547 15962 18547 0 net24
rlabel metal2 25530 23341 25530 23341 0 net25
rlabel metal2 15686 19244 15686 19244 0 net26
rlabel metal1 24518 12648 24518 12648 0 net27
rlabel metal2 24058 13498 24058 13498 0 net28
rlabel metal1 22908 17170 22908 17170 0 net29
rlabel metal1 9108 17102 9108 17102 0 net3
rlabel metal1 23874 10710 23874 10710 0 net30
rlabel metal1 4140 14042 4140 14042 0 net31
rlabel metal1 11362 10778 11362 10778 0 net32
rlabel metal1 25668 12818 25668 12818 0 net33
rlabel metal1 8602 3060 8602 3060 0 net34
rlabel metal1 7038 19856 7038 19856 0 net35
rlabel metal1 8648 16762 8648 16762 0 net36
rlabel metal1 23092 16762 23092 16762 0 net37
rlabel metal1 22305 16150 22305 16150 0 net38
rlabel via2 12558 13379 12558 13379 0 net39
rlabel metal2 3726 14280 3726 14280 0 net4
rlabel metal2 7682 15674 7682 15674 0 net40
rlabel metal1 6854 16048 6854 16048 0 net41
rlabel metal1 16606 21964 16606 21964 0 net42
rlabel metal1 13938 23732 13938 23732 0 net43
rlabel metal1 10166 25296 10166 25296 0 net44
rlabel metal2 26450 14518 26450 14518 0 net45
rlabel metal1 10350 4250 10350 4250 0 net46
rlabel metal1 16422 6324 16422 6324 0 net47
rlabel metal1 20240 15538 20240 15538 0 net48
rlabel metal2 7222 14212 7222 14212 0 net49
rlabel metal2 1610 15827 1610 15827 0 net5
rlabel metal2 23966 16371 23966 16371 0 net50
rlabel metal2 19274 8466 19274 8466 0 net51
rlabel metal2 14122 4386 14122 4386 0 net52
rlabel metal2 13018 24888 13018 24888 0 net53
rlabel metal1 14904 26282 14904 26282 0 net54
rlabel metal1 6486 26962 6486 26962 0 net55
rlabel metal2 9706 14212 9706 14212 0 net56
rlabel metal2 19090 15164 19090 15164 0 net57
rlabel metal2 21942 23902 21942 23902 0 net58
rlabel metal1 4922 4182 4922 4182 0 net59
rlabel metal2 1610 17408 1610 17408 0 net6
rlabel metal1 19366 12886 19366 12886 0 net60
rlabel metal1 4830 20570 4830 20570 0 net61
rlabel metal1 25116 14994 25116 14994 0 net62
rlabel metal1 6348 14994 6348 14994 0 net63
rlabel metal2 14306 16320 14306 16320 0 net64
rlabel metal1 4416 7514 4416 7514 0 net65
rlabel metal1 4370 15470 4370 15470 0 net66
rlabel metal2 14122 14144 14122 14144 0 net67
rlabel metal1 19136 6766 19136 6766 0 net68
rlabel metal2 6394 3196 6394 3196 0 net69
rlabel metal2 1610 19737 1610 19737 0 net7
rlabel metal2 1610 20893 1610 20893 0 net8
rlabel metal1 26082 8942 26082 8942 0 net9
<< properties >>
string FIXED_BBOX 0 0 27988 30132
<< end >>
