* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt level_shifter level_shifter_0/VDD level_shifter_0/VH level_shifter_0/GND level_shifter_0/IN
+ level_shifter_0/OUT
X0 a_1660_2346# level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X2 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X3 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X4 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X5 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X6 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X7 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X8 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X9 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X10 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X11 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X12 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X13 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.6 as=2.9 ps=20.3 w=20 l=0.5
X14 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X15 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X16 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X17 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X18 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X19 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X20 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X21 level_shifter_0/cruzados_0/OUT level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X22 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X23 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X24 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X25 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X26 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X27 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X28 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X29 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X30 level_shifter_0/VDD level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X31 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X32 level_shifter_0/cruzados_0/OUT a_1660_2346# level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X33 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X34 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=5.8 ps=40.6 w=20 l=0.5
X35 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X36 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X37 level_shifter_0/cruzados_0/OUT level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X38 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X39 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X40 level_shifter_0/GND level_shifter_0/IN a_1660_2346# level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X41 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X42 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=5.8 ps=40.6 w=20 l=0.5
X43 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X44 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X45 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X46 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X47 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X48 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X49 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X50 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X51 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X52 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X53 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X54 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X55 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X56 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X57 level_shifter_0/GND level_shifter_0/inv_1_8_0/OUT level_shifter_0/cruzados_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X58 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X59 a_1660_2346# level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X60 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=5.8 pd=40.6 as=2.9 ps=20.3 w=20 l=0.5
X61 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X62 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X63 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X64 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X65 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X66 level_shifter_0/VDD level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X67 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X68 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X69 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X70 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X71 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X72 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X73 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X74 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X75 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X76 a_1660_2346# level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X77 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
.ends

.subckt nmos_drain_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# a_100_62#
+ m5_788_894# m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.78 ps=18.8 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.78 pd=18.8 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.86 ps=16.6 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=6.86 pd=16.6 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_lt m4_n1950_0# m4_648_1020# m5_n1950_0# a_n950_0# m5_788_894#
+ m3_n1950_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_n950_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=12.5 ps=32.6 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020# a_1550_0#
X0 a_162_1100# a_0_0# a_100_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.03 ps=14.1 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.1 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.23 ps=16.3 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=6.23 pd=16.3 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_lt m4_648_1020# m3_n950_0# a_n950_0# m4_n950_0# m5_n950_0#
+ m5_788_894# a_0_0# a_162_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_162_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=4.05 ps=28.2 w=4.38 l=0.5
.ends

.subckt nmos_waffle_36x36 dw_n6950_n7050# a_n938_0# a_37562_0# a_n1100_n1200#
Xnmos_drain_in_530 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_541 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_552 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_563 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_574 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_360 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_371 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_382 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_393 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_190 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_509 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_520 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_531 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_542 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_553 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_564 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_575 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_350 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_361 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_372 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_383 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_394 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_180 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_191 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_510 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_521 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_532 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_543 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_554 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_565 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_576 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_340 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_351 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_362 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_373 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_384 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_395 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_170 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_181 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_192 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_490 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_500 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_511 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_522 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_533 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_544 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_555 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_566 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_577 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_330 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_341 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_352 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_363 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_374 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_385 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_396 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_160 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_171 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_182 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_193 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_491 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_480 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_501 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_512 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_523 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_534 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_545 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_556 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_567 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_320 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_331 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_342 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_353 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_364 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_375 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_386 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_397 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_150 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_161 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_172 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_183 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_30 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_194 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_492 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_481 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_470 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_502 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_513 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_524 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_535 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_546 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_557 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_568 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_0 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_310 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_321 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_332 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_343 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_354 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_365 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_376 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_387 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_398 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_140 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_151 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_162 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_173 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_184 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_195 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_20 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_31 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_482 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_493 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_471 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_460 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_503 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_514 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_525 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_536 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_547 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_558 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_569 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_1 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_300 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_311 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_322 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_333 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_344 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_355 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_366 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_377 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_388 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_399 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_130 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_141 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_152 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_163 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_174 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_185 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_196 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_10 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_21 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_32 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_483 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_494 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_472 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_461 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_450 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_504 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_515 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_526 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_537 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_548 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_559 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_2 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_301 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_312 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_323 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_334 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_345 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_356 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_367 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_378 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_389 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_120 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_131 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_142 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_153 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_164 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_175 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_186 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_197 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_11 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_22 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_33 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_484 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_495 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_473 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_462 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_451 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_505 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_516 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_527 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_538 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_549 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_3 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_302 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_313 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_324 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_335 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_346 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_357 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_368 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_379 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_110 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_121 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_132 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_143 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_154 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_165 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_176 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_187 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_198 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_12 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_23 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_485 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_496 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_474 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_463 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_452 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_506 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_517 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_528 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_539 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_4 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_303 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_314 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_325 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_336 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_347 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_358 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_369 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_100 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_111 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_122 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_133 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_144 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_155 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_166 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_177 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_188 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_13 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_24 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_199 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_486 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_497 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_475 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_464 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_453 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_507 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_518 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_529 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_5 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_304 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_315 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_326 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_337 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_348 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_359 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_101 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_112 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_123 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_134 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_145 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_156 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_167 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_178 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_189 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_14 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_25 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_487 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_498 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_476 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_465 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_454 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_508 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_519 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_0 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_6 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_305 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_316 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_327 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_338 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_349 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_102 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_113 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_124 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_135 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_146 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_157 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_168 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_179 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_15 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_26 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_488 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_499 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_477 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_466 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_455 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_509 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_1 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_7 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_306 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_317 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_328 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_339 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_103 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_114 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_125 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_136 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_147 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_158 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_169 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_16 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_27 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_489 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_478 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_467 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_456 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_90 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_2 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_8 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_307 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_318 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_329 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_104 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_115 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_126 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_137 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_148 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_159 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_17 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_28 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_479 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_468 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_457 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_490 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_0 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_80 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_91 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_9 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_3 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_308 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_319 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_105 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_116 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_127 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_138 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_149 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_18 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_29 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_469 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_458 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_480 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_491 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_1 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_70 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_81 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_92 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_4 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_309 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_106 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_117 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_128 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_139 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_19 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_459 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_470 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_481 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_492 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_2 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_60 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_71 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_82 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_93 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_5 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_107 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_118 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_129 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_460 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_471 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_482 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_493 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_3 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_290 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_50 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_61 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_72 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_83 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_94 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_6 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_108 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_119 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_450 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_461 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_472 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_483 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_494 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_4 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_280 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_291 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_40 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_51 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_62 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_73 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_84 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_95 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_7 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_109 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_440 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_451 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_462 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_473 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_484 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_495 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_5 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_270 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_281 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_292 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_30 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_41 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_52 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_63 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_74 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_85 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_96 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_8 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_430 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_441 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_452 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_463 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_474 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_485 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_496 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_6 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_260 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_271 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_282 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_293 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_20 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_31 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_42 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_53 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_64 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_75 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_86 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_97 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_9 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_420 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_431 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_442 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_453 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_464 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_475 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_486 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_497 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_7 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_250 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_261 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_272 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_283 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_294 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_10 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_21 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_32 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_43 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_54 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_65 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_76 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_87 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_98 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_570 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_30 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_410 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_421 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_432 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_443 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_454 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_465 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_476 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_487 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_498 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_8 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_240 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_251 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_262 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_273 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_284 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_295 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_11 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_22 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_33 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_44 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_55 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_560 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_571 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_66 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_77 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_88 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_99 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_20 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_31 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_400 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_411 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_422 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_433 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_444 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_455 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_466 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_477 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_488 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_499 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_9 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_230 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_241 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_252 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_263 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_274 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_285 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_296 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_30 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_12 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_23 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_34 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_45 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_56 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_67 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_78 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_89 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_550 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_561 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_572 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_10 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_21 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_32 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_401 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_412 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_423 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_434 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_445 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_456 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_467 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_478 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_489 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_220 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_231 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_242 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_253 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_264 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_275 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_286 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_297 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_20 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_31 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_13 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_24 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_35 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_46 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_57 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_68 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_79 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_540 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_551 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_562 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_573 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_11 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_22 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_33 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_0 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_402 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_413 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_424 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_435 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_446 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_457 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_468 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_479 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_10 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_21 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_32 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_210 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_221 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_232 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_243 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_254 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_265 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_276 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_287 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_298 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_14 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_25 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_36 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_47 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_58 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_69 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_530 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_541 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_552 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_563 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_574 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_12 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_23 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_1 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_403 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_414 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_425 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_436 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_447 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_458 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_469 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_200 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_211 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_222 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_233 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_244 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_255 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_266 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_277 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_288 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_299 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_11 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_22 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_33 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_15 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_26 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_37 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_48 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_59 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_520 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_531 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_542 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_553 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_564 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_575 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_13 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_24 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_2 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_404 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_415 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_426 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_437 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_448 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_459 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_201 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_212 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_223 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_234 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_245 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_256 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_267 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_278 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_289 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_12 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_23 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_16 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_27 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_38 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_49 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_510 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_521 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_532 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_543 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_554 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_565 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_576 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_14 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_25 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_3 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_405 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_416 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_427 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_438 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_449 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_202 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_213 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_224 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_235 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_246 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_257 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_268 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_279 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_13 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_24 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_500 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_511 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_522 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_533 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_544 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_555 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_17 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_28 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_39 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_566 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_577 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_15 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_26 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_4 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_406 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_417 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_428 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_439 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_203 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_214 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_225 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_236 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_247 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_258 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_269 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_14 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_25 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_18 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_29 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_501 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_512 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_523 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_534 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_545 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_556 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_567 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_16 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_27 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_5 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_407 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_418 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_429 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_204 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_15 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_26 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_215 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_226 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_237 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_248 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_259 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_19 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_502 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_513 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_524 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_535 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_546 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_557 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_568 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_17 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_28 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_6 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_408 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_419 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_205 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_216 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_227 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_238 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_249 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_16 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_27 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_503 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_514 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_525 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_536 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_547 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_558 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_569 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_18 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_29 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_7 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_409 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_206 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_217 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_228 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_239 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_17 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_28 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_504 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_515 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_526 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_537 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_548 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_559 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_570 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_19 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_8 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_207 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_218 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_229 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_18 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_29 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_505 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_516 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_527 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_538 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_549 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_560 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_571 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_390 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_9 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_208 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_219 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_19 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_506 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_517 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_528 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_539 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_550 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_561 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_572 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_380 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_391 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_209 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_507 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_518 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_529 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_540 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_551 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_562 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_573 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_370 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_381 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_392 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_508 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_519 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
X0 a_37562_0# a_n1100_n1200# a_n938_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X1 a_37562_0# a_n1100_n1200# a_n938_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_n938_0# a_n1100_n1200# a_37562_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_37562_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt power_stage_3 nmos_waffle_36x36_1/dw_n6950_n7050# VP out nmos_waffle_36x36_0/dw_n6950_n7050#
+ s2 s1 VN
Xnmos_waffle_36x36_0 nmos_waffle_36x36_0/dw_n6950_n7050# out VN s1 nmos_waffle_36x36
Xnmos_waffle_36x36_1 nmos_waffle_36x36_1/dw_n6950_n7050# VP out s2 nmos_waffle_36x36
.ends

.subckt mimcap_30x30 c2_30_30# c1_30_30# m3_0_0#
X0 c1_30_30# m3_0_0# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X1 c2_30_30# c1_30_30# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt mimcap_210x420 mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0# mimcap_30x30_9/c2_30_30#
Xmimcap_30x30_90 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_80 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_91 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_70 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_81 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_92 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_60 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_71 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_82 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_93 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_50 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_61 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_72 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_83 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_94 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_40 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_51 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_62 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_73 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_84 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_95 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_96 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_30 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_41 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_52 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_63 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_74 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_85 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_97 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_20 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_31 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_42 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_53 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_64 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_75 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_86 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_21 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_10 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_32 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_43 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_54 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_65 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_76 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_87 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_22 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_11 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_0 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_33 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_44 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_55 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_66 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_77 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_88 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_23 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_12 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_34 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_45 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_56 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_67 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_78 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_89 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_1 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_2 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_24 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_13 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_35 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_46 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_57 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_68 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_79 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_14 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_25 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_36 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_47 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_58 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_69 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_3 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_15 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_4 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_26 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_37 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_48 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_59 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_16 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_27 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_38 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_49 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_5 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_17 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_28 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_39 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_6 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_18 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_29 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_7 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_19 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_8 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_9 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
.ends

.subckt bootstrap_diode a_138_138# dw_n206_n206#
D0 dw_n206_n206# a_138_138# sky130_fd_pr__diode_pw2nd_05v5 pj=5.08e+07 area=1.6129e+14
.ends

.subckt boot_ls_stage w_n1158_n782# VRE Vboot RESET V5v0LS SET VFE GND
X0 V5v0LS a_n824_n1882# GND sky130_fd_pr__res_xhigh_po_0p35 l=2.61
X1 Vboot RESET RESET Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X2 a_n1778_n1384# a_n824_n1218# GND sky130_fd_pr__res_xhigh_po_0p35 l=2.61
X3 w_n1158_n782# a_n824_n1218# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X4 Vboot RESET w_n1370_986# Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 GND a_n824_n1218# w_n1158_n782# GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
X7 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_n1778_n1384# a_n824_n1550# GND sky130_fd_pr__res_xhigh_po_0p35 l=2.61
X9 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 SET SET Vboot Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X12 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 SET SET w_n1370_986# w_n1370_986# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 w_888_986# RESET RESET w_888_986# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 w_888_986# SET Vboot Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 GND a_n824_n1218# a_n824_n1218# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X19 Vboot SET RESET Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=1
X20 a_n1778_n1716# a_n824_n1882# GND sky130_fd_pr__res_xhigh_po_0p35 l=2.61
X21 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X22 SET RESET Vboot Vboot sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=1
X23 a_n1778_n1716# a_n824_n1550# GND sky130_fd_pr__res_xhigh_po_0p35 l=2.61
X24 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X26 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X27 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt buffer QN Vout Q VDD VSS
X0 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X1 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 VSS Q a_n195_154# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X4 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X7 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_n137_16# a_n195_154# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.475 ps=3.37 w=3 l=0.5
X10 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X11 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X12 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X13 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X14 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X16 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X17 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X18 VDD a_n137_16# a_n195_154# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.475 pd=3.37 as=0.29 ps=2.58 w=1 l=0.5
X19 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X20 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X21 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X22 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=3.14 ps=22.3 w=10.8 l=0.5
X23 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X24 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X25 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X26 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=3.14 pd=22.3 as=1.57 ps=11.1 w=10.8 l=0.5
X27 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X28 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X29 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X30 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X31 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X32 a_n137_16# QN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X33 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X34 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X35 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X36 Vout a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X37 Vout a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X38 VDD a_n137_16# Vout VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X39 VSS a_n137_16# Vout VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VPWR X VNB VPB
X0 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.33 as=0.213 ps=2.16 w=0.82 l=0.5
X1 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.217 pd=2.17 as=0.17 ps=1.36 w=0.82 l=0.5
X2 VPWR a_390_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.138 ps=1.27 w=1 l=0.15
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.36 as=0.27 ps=2.54 w=1 l=0.15
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.158 ps=1.33 w=1 l=0.15
X5 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=0.098 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.5
X6 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.01 as=0.113 ps=1.38 w=0.42 l=0.15
X7 VGND a_390_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.164 pd=1.62 as=0.0578 ps=0.695 w=0.42 l=0.15
X8 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=1.01 w=0.65 l=0.5
X9 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.098 ps=0.98 w=0.42 l=0.15
.ends

.subckt sp_delay sky130_fd_sc_hd__clkdlybuf4s50_2_0/A sky130_fd_sc_hd__clkdlybuf4s50_2_5/X
+ sky130_fd_sc_hd__tap_1_1/VPB VSUBS
Xsky130_fd_sc_hd__clkdlybuf4s50_2_0 sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_1/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_1 sky130_fd_sc_hd__clkdlybuf4s50_2_1/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_2/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_2 sky130_fd_sc_hd__clkdlybuf4s50_2_2/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_3/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_3 sky130_fd_sc_hd__clkdlybuf4s50_2_3/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_4/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_4 sky130_fd_sc_hd__clkdlybuf4s50_2_4/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_5/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
Xsky130_fd_sc_hd__clkdlybuf4s50_2_5 sky130_fd_sc_hd__clkdlybuf4s50_2_5/A VSUBS sky130_fd_sc_hd__tap_1_1/VPB
+ sky130_fd_sc_hd__clkdlybuf4s50_2_5/X VSUBS sky130_fd_sc_hd__tap_1_1/VPB sky130_fd_sc_hd__clkdlybuf4s50_2
.ends

.subckt sp_delay2x VIN VOUT VSS VCC
Xsp_delay_0 VIN sp_delay_1/sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VCC VSS sp_delay
Xsp_delay_1 sp_delay_1/sky130_fd_sc_hd__clkdlybuf4s50_2_0/A VOUT VCC VSS sp_delay
.ends

.subckt sp_delay_top VCC VIN VOUT VSS
Xsp_delay2x_0 VIN sp_delay2x_1/VIN VSS VCC sp_delay2x
Xsp_delay2x_1 sp_delay2x_1/VIN sp_delay2x_2/VIN VSS VCC sp_delay2x
Xsp_delay2x_2 sp_delay2x_2/VIN VOUT VSS VCC sp_delay2x
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VPWR X VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt short_pulse_generator Vin VFE VRE VCC VSS
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A VSS VCC sp_delay_top_0/VIN VSS
+ VCC sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_2_0 Vin VSS VCC sky130_fd_sc_hd__inv_2_0/Y VSS VCC sky130_fd_sc_hd__inv_2
Xsp_delay_top_0 VCC sp_delay_top_0/VIN sp_delay_top_0/VOUT VSS sp_delay_top
Xsky130_fd_sc_hd__and2_2_0 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_8_0/A VSS
+ VCC VRE VSS VCC sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__and2_2_1 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/A VSS
+ VCC VFE VSS VCC sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__inv_1_1 sp_delay_top_0/VOUT VSS VCC sky130_fd_sc_hd__inv_1_2/A VSS
+ VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_2_0/Y VSS VCC sky130_fd_sc_hd__inv_8_0/A
+ VSS VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VSS VCC sky130_fd_sc_hd__inv_1_2/Y
+ VSS VCC sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_8_0/A VSS VCC sky130_fd_sc_hd__inv_1_3/Y
+ VSS VCC sky130_fd_sc_hd__inv_1
.ends

.subckt nand_5v NAND B A VDD VSS
X0 a_n29_n1168# B VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
X1 NAND B VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
X2 NAND A a_n29_n1168# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
X3 VDD A NAND VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
.ends

.subckt driver_bootstrap buffer_0/Vout boot_ls_stage_0/V5v0LS w_n3969_322# short_pulse_generator_0/Vin
+ VBOOT VSUBS short_pulse_generator_0/VCC VSource
Xboot_ls_stage_0 w_n3969_322# boot_ls_stage_0/VRE VBOOT nand_5v_1/A boot_ls_stage_0/V5v0LS
+ nand_5v_0/A boot_ls_stage_0/VFE VSUBS boot_ls_stage
Xbuffer_0 nand_5v_1/B buffer_0/Vout buffer_0/Q VBOOT VSource buffer
Xshort_pulse_generator_0 short_pulse_generator_0/Vin boot_ls_stage_0/VFE boot_ls_stage_0/VRE
+ short_pulse_generator_0/VCC VSUBS short_pulse_generator
Xnand_5v_1 buffer_0/Q nand_5v_1/B nand_5v_1/A VBOOT VSource nand_5v
Xnand_5v_0 nand_5v_1/B buffer_0/Q nand_5v_0/A VBOOT VSource nand_5v
.ends

.subckt converter_3 V1v8 driver_bootstrap_0/short_pulse_generator_0/Vin V5v0LS VDD
+ VSS level_shifter_0/level_shifter_0/IN w_113334_n12600# Vout
Xlevel_shifter_0 V1v8 V5v0LS VSS level_shifter_0/level_shifter_0/IN power_stage_3_0/s1
+ level_shifter
Xpower_stage_3_0 VDD VDD Vout VDD power_stage_3_0/s2 power_stage_3_0/s1 VSS power_stage_3
Xmimcap_210x420_0 Vboot Vout Vout mimcap_210x420
Xbootstrap_diode_0 Vboot V5v0LS bootstrap_diode
Xdriver_bootstrap_0 power_stage_3_0/s2 V5v0LS w_113334_n12600# driver_bootstrap_0/short_pulse_generator_0/Vin
+ Vboot VSS V1v8 Vout driver_bootstrap
.ends

.subckt pmos_source_in m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# m5_788_894# m4_0_0#
+ a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.86 ps=16.6 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=6.86 pd=16.6 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_drain_in m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.78 ps=18.8 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=2.78 pd=18.8 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_source_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.23 ps=16.3 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=6.23 pd=16.3 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_source_frame_lt m4_n1950_0# m4_648_1020# w_n1150_0# m5_n1950_0# m5_788_894#
+ m3_n1950_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_n1150_0# w_n1150_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=12.5 ps=32.6 w=4.38 l=0.5
.ends

.subckt pmos_drain_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# w_0_0# a_100_62#
+ m5_788_894# m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.03 ps=14.1 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=2.03 pd=14.1 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt pmos_drain_frame_lt m4_648_1020# w_n1150_0# m3_n950_0# m4_n950_0# m5_n950_0#
+ m5_788_894# a_0_0# a_162_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_162_0# w_n1150_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=4.05 ps=28.2 w=4.38 l=0.5
.ends

.subckt pmos_waffle_48x48 a_n938_0# a_n1100_n1200# a_50762_0#
Xpmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_802 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_813 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_824 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_835 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_846 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_857 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_868 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_879 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_603 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_614 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_625 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_636 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_647 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_658 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_669 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_38 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1051 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1040 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_643 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_632 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_621 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_610 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_676 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_687 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_698 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_665 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_654 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_400 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_411 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_422 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_433 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_444 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_455 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_466 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_477 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_488 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_499 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_495 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_484 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_473 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_462 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_451 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_230 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_241 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_252 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_263 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_274 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_285 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_296 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_29 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_18 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_53 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_64 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_75 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_86 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_97 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1049 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1038 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1027 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1016 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1005 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_829 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_818 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_807 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_803 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_814 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_825 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_836 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_847 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_858 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_869 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_604 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_615 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_626 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_637 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_648 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_659 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_39 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1052 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1041 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1030 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_677 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_666 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_655 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_644 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_633 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_622 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_611 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_600 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_688 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_699 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_401 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_412 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_423 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_434 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_445 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_456 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_467 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_478 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_489 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_990 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_496 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_485 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_474 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_463 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_452 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_220 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_231 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_242 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_253 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_264 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_275 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_286 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_297 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_19 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_54 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_65 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_76 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_87 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_98 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1039 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1028 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1017 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1006 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_819 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_808 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_804 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_815 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_826 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_837 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_848 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_859 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_605 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_616 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_627 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_638 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_649 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1042 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1031 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1020 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1053 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_678 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_689 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_667 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_656 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_645 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_634 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_623 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_612 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_601 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_402 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_413 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_424 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_435 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_446 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_457 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_468 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_479 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_991 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_980 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_497 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_486 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_475 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_464 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_453 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_210 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_221 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_232 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_243 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_254 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_265 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_276 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_287 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_298 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_55 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_66 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_77 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_88 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_99 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1029 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1018 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1007 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_809 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_805 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_816 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_827 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_838 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_849 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_606 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_617 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_628 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_639 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1054 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1043 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1032 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1021 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1010 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_679 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_668 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_657 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_646 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_635 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_624 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_613 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_602 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_403 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_414 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_425 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_436 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_447 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_458 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_469 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_992 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_981 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_970 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_498 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_487 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_476 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_465 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_454 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_200 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_211 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_222 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_233 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_244 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_255 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_266 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_277 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_288 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_299 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_56 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_67 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_78 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_89 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1019 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1008 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_806 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_817 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_828 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_839 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_607 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_618 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_629 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1055 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1044 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1033 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1022 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1011 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1000 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_625 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_614 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_603 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_669 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_658 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_647 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_636 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_404 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_415 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_426 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_437 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_448 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_459 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_993 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_982 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_971 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_960 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_477 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_466 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_455 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_499 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_488 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_201 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_212 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_223 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_234 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_245 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_256 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_267 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_278 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_289 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_790 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_46 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_57 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_68 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_79 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1009 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_807 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_818 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_829 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_608 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_619 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1056 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1045 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1034 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1023 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1012 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1001 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_659 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_648 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_637 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_626 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_615 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_604 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_405 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_416 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_427 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_438 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_449 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_994 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_983 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_972 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_961 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_950 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_489 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_478 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_467 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_456 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_202 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_213 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_224 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_235 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_246 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_257 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_268 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_279 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_990 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_791 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_780 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_47 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_58 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_69 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_808 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_819 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_609 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1024 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1013 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1002 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1057 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1046 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1035 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_649 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_638 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_627 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_616 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_605 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_406 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_417 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_428 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_439 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_951 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_940 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_995 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_984 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_973 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_962 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_479 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_468 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_457 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_203 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_214 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_225 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_236 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_247 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_258 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_269 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_991 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_980 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_792 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_781 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_770 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_48 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_59 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_809 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1047 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1036 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1025 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1014 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1003 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_639 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_628 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_617 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_606 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_407 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_418 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_429 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_985 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_974 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_963 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_952 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_941 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_930 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_996 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_469 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_458 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_204 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_215 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_226 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_237 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_248 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_259 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_981 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_970 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_992 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_793 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_782 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_771 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_760 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_590 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_49 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1048 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1037 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1026 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1015 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1004 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_607 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_629 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_618 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_408 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_419 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_997 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_986 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_975 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_964 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_953 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_942 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_931 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_920 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_459 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_205 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_216 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_227 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_238 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_249 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_960 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_993 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_982 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_971 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_794 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_783 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_772 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_761 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_750 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_790 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_580 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_591 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1049 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1038 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1027 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1016 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1005 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_619 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_608 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_409 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_998 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_987 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_976 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_965 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_954 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_943 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_932 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_921 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_910 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_206 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_217 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_228 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_239 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_950 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_961 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_994 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_983 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_972 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_740 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_795 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_784 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_773 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_762 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_751 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_780 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_791 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_570 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_581 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_592 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1006 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1039 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1028 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1017 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_609 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_933 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_922 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_911 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_900 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_999 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_988 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_977 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_966 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_955 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_944 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_207 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_218 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_229 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_940 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_951 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_995 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_984 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_973 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_962 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_774 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_763 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_752 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_741 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_730 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_796 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_785 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_770 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_781 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_792 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_560 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_571 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_582 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_593 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_390 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1029 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1018 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1007 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_967 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_956 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_945 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_934 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_923 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_912 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_901 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_989 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_978 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_208 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_219 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_930 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_941 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_952 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_963 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_996 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_985 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_974 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_797 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_786 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_775 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_764 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_753 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_742 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_731 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_720 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_760 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_771 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_782 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_793 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_550 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_561 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_572 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_583 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_594 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_590 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_380 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_391 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1019 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_1008 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_979 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_968 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_957 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_946 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_935 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_924 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_913 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_902 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_209 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_920 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_931 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_942 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_953 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_997 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_986 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_975 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_964 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_798 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_787 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_776 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_765 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_754 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_743 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_732 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_721 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_710 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_750 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_761 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_772 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_783 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_794 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_540 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_551 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_562 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_573 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_584 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_595 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_591 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_580 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_370 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_381 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_392 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_1009 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_969 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_958 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_947 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_936 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_925 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_914 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_903 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_910 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_921 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_932 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_943 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_954 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_998 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_987 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_976 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_965 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_722 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_711 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_700 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_799 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_788 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_777 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_766 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_755 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_744 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_733 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_740 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_751 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_762 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_773 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_784 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_795 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_530 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_541 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_552 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_563 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_574 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_585 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_596 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_570 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_592 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_581 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_360 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_371 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_382 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_393 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_190 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_915 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_904 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_959 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_948 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_937 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_926 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_900 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_911 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_922 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_933 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_944 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_955 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_999 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_988 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_977 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_966 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_756 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_745 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_734 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_723 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_712 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_701 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_789 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_778 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_767 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_730 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_741 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_752 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_763 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_774 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_785 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_796 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_520 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_531 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_542 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_553 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_564 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_575 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_586 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_597 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_593 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_582 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_571 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_560 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_350 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_361 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_372 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_383 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_394 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_180 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_191 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_949 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_938 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_927 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_916 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_905 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_901 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_912 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_923 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_934 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_945 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_956 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_989 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_978 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_967 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_779 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_768 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_757 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_746 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_735 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_724 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_713 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_702 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_720 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_731 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_742 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_753 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_764 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_775 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_786 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_797 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_510 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_521 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_532 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_543 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_554 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_565 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_576 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_587 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_598 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_594 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_583 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_572 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_561 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_550 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_340 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_351 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_362 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_373 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_384 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_395 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_170 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_181 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_192 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_939 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_928 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_917 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_906 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_902 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_913 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_924 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_935 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_946 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_957 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_968 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_979 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_769 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_758 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_747 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_736 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_725 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_714 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_703 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_710 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_721 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_732 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_743 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_754 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_765 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_776 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_787 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_798 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_500 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_511 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_522 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_533 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_544 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_555 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_566 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_577 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_588 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_599 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_595 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_584 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_573 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_562 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_551 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_540 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_330 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_341 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_352 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_363 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_374 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_385 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_396 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_160 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_171 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_182 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_193 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_929 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_918 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_907 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_903 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_914 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_925 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_936 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_947 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_958 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_969 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_704 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_759 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_748 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_737 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_726 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_715 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_700 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_711 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_722 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_733 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_744 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_755 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_766 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_777 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_788 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_799 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_501 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_512 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_523 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_534 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_545 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_556 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_567 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_578 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_589 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_552 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_541 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_530 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_596 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_585 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_574 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_563 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_320 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_331 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_342 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_353 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_364 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_375 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_386 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_397 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_150 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_161 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_172 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_183 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_194 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_919 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_908 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_904 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_915 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_926 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_937 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_948 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_959 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_738 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_727 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_716 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_705 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_749 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_701 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_712 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_723 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_734 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_745 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_756 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_767 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_778 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_789 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_502 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_513 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_524 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_535 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_546 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_557 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_568 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_579 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_586 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_575 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_564 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_553 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_542 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_531 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_520 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_597 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_310 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_321 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_332 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_343 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_354 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_365 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_376 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_387 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_398 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_140 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_151 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_162 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_173 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_184 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_195 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_909 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_905 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_916 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_927 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_938 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_949 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_739 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_728 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_717 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_706 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_702 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_713 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_724 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_735 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_746 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_757 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_768 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_779 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_503 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_514 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_525 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_536 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_547 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_558 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_569 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_598 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_587 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_576 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_565 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_554 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_543 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_532 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_521 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_510 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_300 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_311 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_322 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_333 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_344 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_355 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_366 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_377 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_388 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_399 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_130 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_141 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_152 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_163 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_174 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_185 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_196 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_906 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_917 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_928 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_939 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_729 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_718 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_707 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_703 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_714 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_725 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_736 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_747 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_758 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_769 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_504 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_515 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_526 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_537 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_548 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_559 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_500 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_599 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_588 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_577 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_566 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_555 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_544 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_533 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_522 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_511 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_301 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_312 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_323 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_334 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_345 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_356 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_367 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_378 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_389 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_890 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_120 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_131 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_142 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_153 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_164 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_175 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_186 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_197 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_907 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_918 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_929 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_719 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_708 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_704 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_715 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_726 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_737 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_748 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_759 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_505 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_516 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_527 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_538 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_549 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_534 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_523 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_512 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_501 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_589 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_578 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_567 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_556 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_545 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_302 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_313 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_324 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_335 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_346 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_357 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_368 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_379 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_891 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_880 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_110 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_121 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_132 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_143 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_154 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_165 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_176 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_187 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_198 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_908 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_919 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_709 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_705 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_716 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_727 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_738 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_749 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_506 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_517 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_528 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_539 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_568 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_557 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_546 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_535 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_524 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_513 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_502 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_579 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_303 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_314 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_325 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_336 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_347 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_358 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_369 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_892 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_881 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_870 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_100 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_111 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_122 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_133 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_144 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_155 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_166 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_177 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_188 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_199 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_909 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_706 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_717 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_728 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_739 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_507 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_518 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_529 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_569 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_558 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_547 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_536 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_525 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_514 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_503 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_304 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_315 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_326 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_337 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_348 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_359 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_20 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_860 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_31 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_42 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_893 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_882 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_871 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_101 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_112 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_123 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_134 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_145 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_0 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_156 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_167 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_178 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_189 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_690 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_0 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_707 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_718 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_729 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_508 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_519 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_559 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_548 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_537 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_526 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_515 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_504 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_305 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_316 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_327 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_338 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_349 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_10 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_21 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_32 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_43 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_883 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_872 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_861 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_850 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_894 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_102 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_113 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_124 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_135 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_146 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_157 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_168 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_179 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_1 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_890 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_691 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_680 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_1 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_40 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_708 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_719 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_509 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_516 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_505 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_549 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_538 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_527 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_306 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_317 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_328 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_339 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_11 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_22 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_33 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_44 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_895 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_884 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_873 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_862 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_851 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_840 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_103 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_114 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_125 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_136 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_147 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_158 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_169 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_2 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_880 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_891 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_670 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_692 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_681 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_2 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_41 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_30 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_709 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_539 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_528 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_517 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_506 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_307 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_318 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_329 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1050 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_12 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_23 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_34 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_45 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_896 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_885 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_874 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_863 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_852 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_841 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_830 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_104 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_3 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_115 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_126 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_137 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_148 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_159 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_870 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_881 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_892 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_660 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_671 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_693 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_682 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_40 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_3 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_490 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_42 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_31 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_20 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_529 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_518 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_507 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_308 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_319 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1051 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1040 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_842 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_831 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_820 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_13 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_24 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_35 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_897 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_886 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_875 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_864 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_853 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_105 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_116 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_127 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_4 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_138 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_149 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_860 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_871 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_882 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_893 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_650 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_661 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_683 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_672 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_694 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_41 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_4 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_690 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_480 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_491 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_43 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_32 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_21 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_10 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_519 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_508 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_309 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1052 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1041 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1030 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_14 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_25 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_36 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_865 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_854 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_843 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_832 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_821 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_810 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_898 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_887 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_876 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_106 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_117 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_128 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_139 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_5 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_850 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_861 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_872 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_883 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_894 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_640 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_651 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_662 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_695 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_684 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_673 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_42 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_5 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_680 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_691 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_470 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_481 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_492 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_33 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_22 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_11 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_44 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_90 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_509 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1053 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1042 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1031 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1020 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_15 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_26 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_37 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_899 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_888 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_877 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_866 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_855 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_844 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_833 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_822 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_811 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_800 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_107 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_118 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_129 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_6 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_840 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_851 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_862 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_873 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_884 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_895 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_630 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_641 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_652 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_663 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_696 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_685 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_674 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_43 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_6 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_681 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_692 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_670 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_460 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_471 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_482 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_493 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_290 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_45 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_34 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_23 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_12 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_80 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_91 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1054 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1043 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1032 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1021 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1010 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_16 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_27 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_38 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_889 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_878 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_867 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_856 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_845 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_834 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_823 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_812 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_801 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_7 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_108 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_119 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_830 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_841 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_852 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_863 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_874 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_885 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_896 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_620 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_631 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_642 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_653 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_664 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_697 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_686 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_675 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_44 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_7 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_682 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_693 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_671 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_660 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_450 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_461 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_472 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_483 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_494 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_490 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_280 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_291 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_35 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_24 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_13 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_70 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_81 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_92 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1033 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1022 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1011 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1000 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1055 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1044 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_824 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_813 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_802 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_17 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_28 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_39 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_879 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_868 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_857 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_846 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_835 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_109 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_lt_8 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_drain_in_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_820 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_831 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_842 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_853 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_864 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_875 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_886 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_897 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_610 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_621 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_632 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_643 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_654 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_665 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_698 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_687 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_676 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_45 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_34 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_8 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_661 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_650 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_683 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_694 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_672 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_440 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_451 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_462 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_473 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_484 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_495 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_491 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_480 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_270 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_281 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_292 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_36 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_25 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_14 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_60 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_71 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_82 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_93 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1056 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1045 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1034 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1023 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1012 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1001 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_18 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_847 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_836 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_825 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_814 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_803 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_frame_rb_29 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_869 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_858 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_9 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0#
+ a_n1100_n1200# a_n938_0# a_50762_0# a_50762_0# pmos_drain_frame_lt
Xpmos_source_in_810 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_821 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_832 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_843 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_854 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_865 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_876 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_887 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_898 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_600 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_611 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_622 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_633 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_644 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_655 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_666 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_699 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_688 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_677 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_35 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_9 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_684 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_695 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_673 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_662 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_651 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_640 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_430 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_441 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_452 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_463 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_474 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_485 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_496 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_492 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_481 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_470 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_260 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_271 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_282 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_293 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_15 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_37 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_26 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_50 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_61 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_72 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_83 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_94 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1057 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1046 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1035 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1024 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1013 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1002 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_19 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_frame_rb
Xpmos_drain_in_859 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_848 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_837 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_826 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_815 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_804 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_800 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_811 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_822 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_833 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_844 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_855 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_866 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_877 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_888 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_899 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_601 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_612 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_623 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_634 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_645 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_656 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_667 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_689 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_678 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_36 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_674 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_685 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_696 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_663 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_652 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_641 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_630 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_420 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_431 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_442 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_453 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_464 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_475 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_486 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_497 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_493 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_482 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_471 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_460 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_250 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_261 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_272 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_283 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_294 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_38 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_27 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_16 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_40 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_51 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_62 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_73 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_84 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_95 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1047 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1036 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1025 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1014 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1003 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_849 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_838 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_827 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_816 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_805 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_801 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_812 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_823 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_834 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_845 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_856 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_867 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_878 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_889 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_602 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_613 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_624 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_635 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_646 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_657 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_668 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_679 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_37 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_1050 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_675 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_686 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_697 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_664 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_653 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_642 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_631 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_620 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_410 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_421 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_432 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_443 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_454 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_465 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_476 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_487 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_498 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_461 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_450 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_494 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_483 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_472 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_240 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_251 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_262 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_273 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_284 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_295 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_frame_lt_39 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_28 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_17 a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_30 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_41 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_52 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_63 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_74 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_85 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_96 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_source_in_1015 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1004 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1048 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1037 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_1026 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_50762_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_806 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_839 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_828 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
Xpmos_drain_in_817 a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_50762_0# a_n938_0#
+ a_50762_0# a_50762_0# a_n1100_n1200# a_50762_0# a_50762_0# pmos_drain_in
X0 a_50762_0# a_n1100_n1200# a_n938_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X1 a_n938_0# a_n1100_n1200# a_50762_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_50762_0# a_n1100_n1200# a_n938_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_50762_0# a_50762_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt nmos_waffle_32x32 dw_n6950_n7050# a_33162_0# a_n938_0# a_n1100_n1200#
Xnmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_360 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_371 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_382 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_393 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_190 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_350 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_361 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_372 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_383 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_394 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_180 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_191 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_340 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_351 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_362 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_373 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_384 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_395 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_170 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_181 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_192 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_330 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_341 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_352 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_363 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_374 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_385 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_396 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_160 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_171 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_182 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_193 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_320 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_331 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_342 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_353 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_364 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_375 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_386 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_397 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_150 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_161 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_172 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_183 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_194 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_0 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_310 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_321 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_332 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_343 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_354 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_365 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_376 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_387 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_398 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_140 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_151 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_162 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_173 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_184 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_195 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_20 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_1 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_300 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_311 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_322 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_333 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_344 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_355 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_366 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_377 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_388 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_399 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_130 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_141 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_152 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_163 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_174 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_185 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_196 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_10 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_21 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_2 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_301 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_312 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_323 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_334 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_345 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_356 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_367 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_378 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_389 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_120 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_131 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_142 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_153 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_164 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_175 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_186 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_197 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_11 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_22 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_3 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_302 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_313 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_324 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_335 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_346 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_357 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_368 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_379 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_110 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_121 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_132 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_143 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_154 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_165 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_176 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_187 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_198 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_12 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_23 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_4 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_303 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_314 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_325 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_336 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_347 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_358 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_369 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_100 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_111 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_122 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_133 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_144 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_155 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_166 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_177 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_188 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_13 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_24 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_199 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_5 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_304 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_315 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_326 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_337 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_348 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_359 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_101 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_112 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_123 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_134 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_145 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_156 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_167 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_178 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_189 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_14 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_25 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_0 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_6 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_305 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_316 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_327 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_338 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_349 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_102 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_113 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_124 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_135 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_146 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_157 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_168 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_179 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_15 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_26 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_1 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_7 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_306 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_317 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_328 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_339 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_103 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_114 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_125 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_136 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_147 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_158 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_169 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_16 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_27 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_90 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_2 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_8 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_307 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_318 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_329 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_104 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_115 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_126 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_137 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_148 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_159 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_17 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_28 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_0 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_80 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_91 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_9 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_3 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_308 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_319 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_105 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_116 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_127 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_138 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_149 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_18 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_29 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_1 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_70 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_81 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_92 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_4 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_309 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_106 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_117 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_128 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_139 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_19 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_2 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_60 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_71 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_82 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_93 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_5 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_107 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_118 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_129 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_3 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_290 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_50 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_61 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_72 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_83 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_94 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_6 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_in_108 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_119 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_4 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_280 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_291 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_40 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_51 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_62 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_73 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_84 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_95 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_7 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_109 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_440 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_5 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_270 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_281 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_292 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_30 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_41 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_52 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_63 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_74 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_85 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_96 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_8 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_430 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_441 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_6 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_260 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_271 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_282 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_293 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_20 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_31 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_42 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_53 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_64 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_75 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_86 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_97 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_lt_9 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_420 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_431 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_442 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_7 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_250 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_261 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_272 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_283 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_294 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_10 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_21 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_32 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_43 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_54 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_65 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_76 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_87 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_98 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_410 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_421 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_432 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_443 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_8 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_240 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_251 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_262 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_273 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_284 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_295 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_11 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_22 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_33 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_44 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_55 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_66 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_77 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_88 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_99 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_20 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_400 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_411 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_422 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_433 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_444 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_9 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_230 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_241 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_252 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_263 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_274 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_285 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_296 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_12 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_23 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_34 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_45 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_56 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_67 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_78 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_89 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_10 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_21 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_401 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_412 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_423 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_434 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_445 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_220 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_231 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_242 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_253 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_264 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_275 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_286 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_297 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_20 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_13 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_24 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_35 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_46 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_57 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_68 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_79 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_11 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_22 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_0 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_402 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_413 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_424 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_435 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_446 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_10 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_21 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_210 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_221 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_232 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_243 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_254 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_265 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_276 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_287 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_298 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_14 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_25 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_36 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_47 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_58 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_69 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_12 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_23 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_1 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_403 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_414 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_425 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_436 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_447 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_200 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_211 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_222 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_233 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_244 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_255 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_266 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_277 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_288 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_299 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_11 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_22 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_15 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_26 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_37 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_48 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_59 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_13 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_24 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_2 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_404 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_415 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_426 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_437 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_448 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_201 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_212 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_223 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_234 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_245 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_256 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_267 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_278 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_289 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_12 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_23 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_16 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_27 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_38 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_49 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_14 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_25 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_3 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_405 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_416 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_427 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_438 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_449 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_202 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_213 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_224 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_235 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_246 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_257 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_268 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_279 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_13 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_24 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_17 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_28 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_39 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_15 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_26 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_4 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_406 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_417 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_428 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_439 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_203 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_214 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_225 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_236 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_247 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_258 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_269 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_14 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_25 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_18 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_29 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_16 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_27 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_5 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_407 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_418 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_429 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_204 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_15 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_26 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_in_215 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_226 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_237 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_248 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_259 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_19 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_17 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_28 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_6 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_408 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_419 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_205 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_216 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_227 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_238 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_249 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_16 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_27 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_18 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_29 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_7 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_409 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_206 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_217 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_228 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_239 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_17 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_28 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_19 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_33162_0#
+ a_n1100_n1200# a_n938_0# a_33162_0# a_33162_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_8 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_207 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_218 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_229 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_18 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_29 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_390 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_frame_lt_9 a_n938_0# a_n938_0# a_n938_0# a_33162_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_208 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_219 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_frame_rb_19 a_33162_0# a_33162_0# a_33162_0# a_33162_0# a_n938_0# a_33162_0#
+ a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# a_33162_0# nmos_drain_frame_rb
Xnmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_380 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_391 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_209 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_370 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_381 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_drain_in_392 a_33162_0# a_33162_0# a_33162_0# dw_n6950_n7050# a_33162_0# a_33162_0#
+ a_n938_0# a_33162_0# a_33162_0# a_n1100_n1200# a_33162_0# a_33162_0# nmos_drain_in
Xnmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_33162_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
X0 a_n938_0# a_n1100_n1200# a_33162_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X1 a_33162_0# a_n1100_n1200# a_n938_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_33162_0# a_n1100_n1200# a_n938_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_33162_0# a_33162_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt power_stage_1 nmos_waffle_32x32_0/dw_n6950_n7050# out s4 s3 s2 VN s1 VSUBS
+ fc1 fc2 nmos_waffle_32x32_1/dw_n6950_n7050# VP
Xpmos_waffle_48x48_0 out s2 fc1 pmos_waffle_48x48
Xpmos_waffle_48x48_1 fc1 s1 VP pmos_waffle_48x48
Xnmos_waffle_32x32_0 nmos_waffle_32x32_0/dw_n6950_n7050# VN fc2 s4 nmos_waffle_32x32
Xnmos_waffle_32x32_1 nmos_waffle_32x32_1/dw_n6950_n7050# fc2 out s3 nmos_waffle_32x32
.ends

.subckt converter_1 power_stage_1_0/nmos_waffle_32x32_1/dw_n6950_n7050# power_stage_1_0/nmos_waffle_32x32_0/dw_n6950_n7050#
+ D4 D2 D3 VLS m1_2000_83200# power_stage_1_0/fc1 power_stage_1_0/VP power_stage_1_0/VN
+ VDD D1 VSUBS power_stage_1_0/fc2 power_stage_1_0/out
Xlevel_shifter_0 VDD VLS VSUBS D1 power_stage_1_0/s1 level_shifter
Xlevel_shifter_1 VDD VLS VSUBS D2 power_stage_1_0/s2 level_shifter
Xlevel_shifter_2 VDD VLS VSUBS D3 power_stage_1_0/s3 level_shifter
Xlevel_shifter_3 VDD VLS VSUBS D4 power_stage_1_0/s4 level_shifter
Xpower_stage_1_0 power_stage_1_0/nmos_waffle_32x32_0/dw_n6950_n7050# power_stage_1_0/out
+ power_stage_1_0/s4 power_stage_1_0/s3 power_stage_1_0/s2 power_stage_1_0/VN power_stage_1_0/s1
+ VSUBS power_stage_1_0/fc1 power_stage_1_0/fc2 power_stage_1_0/nmos_waffle_32x32_1/dw_n6950_n7050#
+ power_stage_1_0/VP power_stage_1
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VPWR X VNB VPB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VPWR Y VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.223 pd=2.21 as=0.121 ps=1.16 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.121 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VPWR X VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VPWR X VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VPWR X VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VPWR X VNB VPB
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C VGND VPWR X VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.198 pd=1.39 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.128 ps=1.04 w=0.65 l=0.15
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.198 ps=1.39 w=1 l=0.15
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.177 ps=1.36 w=1 l=0.15
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138 ps=1.08 w=0.65 l=0.15
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VPWR X VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VPWR Q VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VPWR X VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VPWR Y VNB VPB
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VPWR X VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VPWR X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VPWR X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VPWR Y VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VPWR X VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VPWR X VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VPWR X VNB VPB
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.109 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.275 ps=1.5 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VPWR X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VPWR X VNB VPB
X0 a_244_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.217 pd=2.17 as=0.193 ps=1.41 w=0.82 l=0.25
X1 VPWR a_244_47# a_355_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.273 pd=1.61 as=0.217 ps=2.17 w=0.82 l=0.25
X2 X a_355_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.273 ps=1.61 w=1 l=0.15
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.41 as=0.27 ps=2.54 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.07 as=0.113 ps=1.38 w=0.42 l=0.15
X5 VGND a_244_47# a_355_47# VNB sky130_fd_pr__nfet_01v8 ad=0.186 pd=1.26 as=0.172 ps=1.83 w=0.65 l=0.25
X6 X a_355_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.83 as=0.186 ps=1.26 w=0.42 l=0.15
X7 a_244_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.07 w=0.65 l=0.25
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VPWR X VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.263 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.213 ps=1.42 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VPWR X VNB VPB
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VPWR X VNB VPB
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0852 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.269 pd=2.12 as=0.0921 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0921 pd=0.99 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0852 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0901 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0901 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.151 ps=1.28 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151 pd=1.28 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt modulator CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT d1[0]
+ d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[5] d2[4] VPWR VGND
XFILLER_0_23_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1270_ _0626_ _0627_ _0512_ VGND VPWR _0628_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0985_ Shift_Register_Inst.data_out\[11\] _0429_ net23 _0441_ VGND VPWR _0442_ VGND
+ VPWR sky130_fd_sc_hd__a31o_4
XFILLER_0_1_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0770_ Signal_Generator_1_90phase_inst.direction _0279_ _0280_ _0263_ _0281_ VGND
+ VPWR _0025_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_1253_ _0513_ _0616_ _0617_ VGND VPWR _0170_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1322_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0009_ _0095_ VGND VPWR Signal_Generator_1_180phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1184_ _0529_ _0558_ _0559_ _0560_ VGND VPWR _0561_ VGND VPWR sky130_fd_sc_hd__a22oi_4
X_0968_ _0419_ _0424_ VGND VPWR _0427_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_46_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0899_ Signal_Generator_2_180phase_inst.count\[2\] _0371_ VGND VPWR _0378_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0822_ _0319_ _0320_ _0310_ VGND VPWR _0321_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0684_ _0182_ _0216_ _0217_ VGND VPWR _0218_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0753_ Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[0\]
+ VGND VPWR _0268_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_3_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1305_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0006_ _0078_ VGND VPWR Signal_Generator_1_0phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1236_ _0603_ VGND VPWR _0167_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1098_ _0515_ VGND VPWR _0093_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1167_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR _0544_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_19_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1021_ _0452_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[2\]
+ _0451_ VGND VPWR _0455_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0805_ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR _0308_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0667_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ _0195_ VGND VPWR _0205_ VGND VPWR sky130_fd_sc_hd__or3_1
X_0736_ _0254_ _0255_ _0245_ VGND VPWR _0256_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_24_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1219_ _0587_ net39 VGND VPWR _0590_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_30_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold30 Signal_Generator_1_180phase_inst.direction VGND VPWR net55 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 Dead_Time_Generator_inst_2.count_dt\[2\] VGND VPWR net66 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1004_ _0449_ VGND VPWR _0066_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0719_ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VPWR _0243_ VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput20 net20 VGND VPWR PMOS1_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0984_ _0439_ Shift_Register_Inst.data_out\[12\] clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR _0441_ VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_0_13_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1252_ net37 net29 VGND VPWR _0617_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1321_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0008_ _0094_ VGND VPWR Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1183_ _0535_ _0541_ _0554_ VGND VPWR _0560_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_46_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0967_ _0426_ VGND VPWR net22 VGND VPWR sky130_fd_sc_hd__buf_1
X_0898_ Signal_Generator_2_180phase_inst.count\[2\] _0374_ VGND VPWR _0377_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0821_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR _0320_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0752_ _0263_ _0267_ VGND VPWR _0027_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0683_ _0187_ _0205_ Shift_Register_Inst.shift_state\[3\] VGND VPWR _0217_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_3_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1235_ _0601_ _0602_ _0561_ VGND VPWR _0603_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1166_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] VGND VPWR
+ _0543_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1304_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0157_ VGND VPWR Dead_Time_Generator_inst_4.go
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1097_ _0515_ VGND VPWR _0092_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1020_ _0452_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0453_ VGND VPWR _0454_ VGND VPWR sky130_fd_sc_hd__o211a_1
X_0804_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0305_ _0306_ VGND VPWR _0307_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0735_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR _0255_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0666_ _0204_ VGND VPWR _0149_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1149_ Shift_Register_Inst.data_out\[16\] net7 VGND VPWR _0526_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_1218_ _0584_ _0586_ _0588_ VGND VPWR _0589_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_27_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold20 Dead_Time_Generator_inst_3.count_dt\[3\] VGND VPWR net45 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 Dead_Time_Generator_inst_1.count_dt\[0\] VGND VPWR net56 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 Shift_Register_Inst.data_out\[17\] VGND VPWR net67 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1003_ _0446_ VGND VPWR _0449_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_16_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0718_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0240_ _0241_ VGND VPWR _0242_ VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_12_110 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0649_ _0189_ _0192_ VGND VPWR _0193_ VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput21 net21 VGND VPWR PMOS1_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0983_ net18 _0432_ _0438_ _0439_ VGND VPWR _0440_ VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_0_22_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1320_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0007_ _0093_ VGND VPWR Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1182_ _0539_ _0540_ _0557_ _0528_ VGND VPWR _0559_ VGND VPWR sky130_fd_sc_hd__a211oi_2
X_1251_ Dead_Time_Generator_inst_3.count_dt\[0\] _0615_ VGND VPWR _0616_ VGND VPWR
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0966_ _0416_ _0417_ _0424_ VGND VPWR _0426_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0897_ _0041_ _0375_ _0376_ VGND VPWR _0036_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0820_ _0309_ VGND VPWR _0319_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0751_ net53 Signal_Generator_1_90phase_inst.count\[4\] _0266_ VGND VPWR _0267_ VGND
+ VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_3_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1303_ clknet_1_1__leaf_CLK_SR _0156_ _0077_ VGND VPWR Shift_Register_Inst.shift_state\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0682_ Shift_Register_Inst.data_out\[8\] VGND VPWR _0216_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1096_ _0515_ VGND VPWR _0091_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1165_ Shift_Register_Inst.data_out\[13\] net6 VGND VPWR _0542_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_1234_ Dead_Time_Generator_inst_2.count_dt\[2\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ _0594_ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VPWR _0602_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0949_ Dead_Time_Generator_inst_4.go net5 _0228_ VGND VPWR _0414_ VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_33_130 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0665_ _0182_ Dead_Time_Generator_inst_1.dt\[3\] _0203_ VGND VPWR _0204_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0803_ Signal_Generator_1_270phase_inst.direction VGND VPWR _0306_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0734_ _0244_ VGND VPWR _0254_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_24_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1217_ _0585_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0587_ VGND VPWR _0588_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1148_ _0519_ _0524_ VGND VPWR _0525_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1079_ _0512_ VGND VPWR _0513_ VGND VPWR sky130_fd_sc_hd__buf_2
Xhold10 Signal_Generator_1_270phase_inst.count\[0\] VGND VPWR net35 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 Signal_Generator_2_90phase_inst.count\[0\] VGND VPWR net46 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 Shift_Register_Inst.shift_state\[1\] VGND VPWR net57 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 Signal_Generator_2_180phase_inst.direction VGND VPWR net68 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1002_ _0448_ VGND VPWR _0065_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0717_ Signal_Generator_1_0phase_inst.direction VGND VPWR _0241_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0648_ _0187_ _0188_ VGND VPWR _0192_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_35_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VPWR PMOS2_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0982_ Shift_Register_Inst.data_out\[11\] VGND VPWR _0439_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_13_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1181_ _0555_ _0556_ _0557_ VGND VPWR _0558_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_1250_ _0611_ _0612_ _0613_ net28 VGND VPWR _0615_ VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_24_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0896_ _0370_ _0375_ net51 VGND VPWR _0376_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0965_ _0425_ VGND VPWR net15 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_40_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1379_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0176_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_0750_ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ _0265_ VGND VPWR _0266_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0681_ _0215_ VGND VPWR _0145_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1233_ Dead_Time_Generator_inst_2.count_dt\[3\] Dead_Time_Generator_inst_2.count_dt\[2\]
+ _0597_ VGND VPWR _0601_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1302_ clknet_1_1__leaf_CLK_SR _0155_ _0076_ VGND VPWR Shift_Register_Inst.shift_state\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1164_ _0228_ _0530_ _0534_ _0539_ _0540_ VGND VPWR _0541_ VGND VPWR sky130_fd_sc_hd__o32a_1
X_1095_ _0515_ VGND VPWR _0090_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0948_ Shift_Register_Inst.data_out\[15\] Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\]
+ VGND VPWR _0413_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_27_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0879_ _0349_ _0360_ _0363_ net52 VGND VPWR _0052_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0802_ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR _0305_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0664_ _0186_ _0187_ _0188_ VGND VPWR _0203_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0733_ _0240_ _0252_ VGND VPWR _0253_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_21_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1216_ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VPWR _0587_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1147_ Signal_Generator_1_0phase_inst.count\[5\] _0520_ _0521_ _0523_ VGND VPWR _0524_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1078_ _0477_ _0494_ _0507_ _0511_ VGND VPWR _0512_ VGND VPWR sky130_fd_sc_hd__o31a_1
Xhold11 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VPWR net36 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 Signal_Generator_2_180phase_inst.count\[0\] VGND VPWR net47 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 Signal_Generator_1_0phase_inst.direction VGND VPWR net58 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 Signal_Generator_2_0phase_inst.direction VGND VPWR net69 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1001_ _0448_ VGND VPWR _0064_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0716_ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VPWR _0240_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0647_ _0190_ _0191_ VGND VPWR _0155_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_35_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput23 net23 VGND VPWR PMOS2_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0981_ net21 _0430_ _0437_ VGND VPWR _0438_ VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_1_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1180_ _0526_ _0527_ _0525_ VGND VPWR _0557_ VGND VPWR sky130_fd_sc_hd__o21ai_1
X_0964_ _0414_ _0424_ VGND VPWR _0425_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_40_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0895_ _0374_ _0371_ VGND VPWR _0375_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_10_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1378_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0175_ VGND VPWR Dead_Time_Generator_inst_2.go
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0680_ _0182_ _0214_ _0190_ VGND VPWR _0215_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1232_ _0581_ _0600_ VGND VPWR _0166_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1301_ clknet_1_1__leaf_CLK_SR _0154_ _0075_ VGND VPWR Shift_Register_Inst.shift_state\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1094_ _0515_ VGND VPWR _0089_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1163_ _0228_ net3 VGND VPWR _0540_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_0947_ _0412_ VGND VPWR net24 VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_27_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0878_ _0361_ _0362_ _0352_ VGND VPWR _0363_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0801_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0287_ _0304_ VGND VPWR _0012_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_24_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0732_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR _0252_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0663_ _0202_ VGND VPWR _0150_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1215_ _0582_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[2\]
+ _0585_ VGND VPWR _0586_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_1146_ _0208_ _0211_ Signal_Generator_1_270phase_inst.count\[5\] _0522_ VGND VPWR
+ _0523_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_46_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1077_ _0477_ _0510_ _0475_ _0476_ VGND VPWR _0511_ VGND VPWR sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold12 Dead_Time_Generator_inst_3.count_dt\[0\] VGND VPWR net37 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 Shift_Register_Inst.shift_state\[4\] VGND VPWR net48 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 Signal_Generator_2_0phase_inst.direction VGND VPWR net59 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1000_ _0448_ VGND VPWR _0063_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0715_ _0239_ VGND VPWR _0135_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0646_ _0186_ _0189_ VGND VPWR _0191_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1129_ _0518_ VGND VPWR _0121_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_35_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VPWR PMOS_PS3 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0980_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] net16
+ VGND VPWR _0437_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_1_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_0963_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] Shift_Register_Inst.data_out\[15\]
+ VGND VPWR _0424_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0894_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ VGND VPWR _0374_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_6_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1377_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0174_ VGND VPWR Dead_Time_Generator_inst_3.count_dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1162_ _0536_ _0537_ _0538_ _0520_ Signal_Generator_1_0phase_inst.count\[0\] VGND
+ VPWR _0539_ VGND VPWR sky130_fd_sc_hd__o32a_1
X_1231_ net66 _0597_ VGND VPWR _0600_ VGND VPWR sky130_fd_sc_hd__xnor2_1
X_1300_ clknet_1_0__leaf_CLK_SR _0153_ _0074_ VGND VPWR Shift_Register_Inst.shift_state\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1093_ _0515_ VGND VPWR _0088_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0946_ net7 Shift_Register_Inst.data_out\[16\] VGND VPWR _0412_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_0877_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VPWR _0362_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_27_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0731_ _0242_ _0249_ _0251_ Signal_Generator_1_0phase_inst.direction VGND VPWR _0002_
+ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0800_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0283_ Signal_Generator_1_180phase_inst.count\[5\] VGND VPWR _0304_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0662_ _0182_ Dead_Time_Generator_inst_1.dt\[2\] _0201_ VGND VPWR _0202_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_1214_ Dead_Time_Generator_inst_2.count_dt\[2\] VGND VPWR _0585_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1145_ _0211_ Signal_Generator_1_90phase_inst.count\[5\] _0208_ VGND VPWR _0522_
+ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_46_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1076_ _0508_ _0492_ _0494_ _0509_ VGND VPWR _0510_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_0929_ _0391_ _0398_ _0400_ Signal_Generator_2_270phase_inst.direction VGND VPWR
+ _0044_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_15_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold13 _0170_ VGND VPWR net38 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 Dead_Time_Generator_inst_1.count_dt\[1\] VGND VPWR net49 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 Shift_Register_Inst.shift_state\[0\] VGND VPWR net60 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0714_ net67 net1 _0238_ VGND VPWR _0239_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0645_ _0186_ _0189_ VGND VPWR _0190_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1128_ _0518_ VGND VPWR _0120_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1059_ _0489_ _0490_ _0485_ VGND VPWR _0493_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_174 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VPWR SIGNAL_OUTPUT VGND VPWR sky130_fd_sc_hd__buf_8
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0962_ _0423_ VGND VPWR net21 VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_0893_ net47 VGND VPWR _0035_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_6_217 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1376_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0173_ VGND VPWR Dead_Time_Generator_inst_3.count_dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1092_ _0515_ VGND VPWR _0087_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1161_ _0208_ _0007_ VGND VPWR _0538_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1230_ _0599_ VGND VPWR _0165_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0876_ _0351_ VGND VPWR _0361_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0945_ _0411_ VGND VPWR net19 VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1359_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0046_ _0132_ VGND VPWR Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0661_ Shift_Register_Inst.shift_state\[3\] _0187_ _0200_ VGND VPWR _0201_ VGND VPWR
+ sky130_fd_sc_hd__or3_1
X_0730_ _0245_ _0250_ VGND VPWR _0251_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1213_ _0582_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0583_ VGND VPWR _0584_ VGND VPWR sky130_fd_sc_hd__o211a_1
X_1144_ _0211_ _0300_ _0208_ VGND VPWR _0521_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1075_ _0503_ _0504_ _0506_ VGND VPWR _0509_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0859_ Signal_Generator_2_90phase_inst.direction VGND VPWR _0348_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0928_ _0394_ _0399_ VGND VPWR _0400_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_30_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold14 Dead_Time_Generator_inst_1.dt\[3\] VGND VPWR net39 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 Dead_Time_Generator_inst_3.count_dt\[1\] VGND VPWR net50 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 Signal_Generator_1_270phase_inst.direction VGND VPWR net61 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0644_ _0187_ _0188_ VGND VPWR _0189_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0713_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ _0237_ VGND VPWR _0238_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_12_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1127_ _0518_ VGND VPWR _0119_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1058_ _0482_ _0483_ _0478_ VGND VPWR _0492_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput15 net15 VGND VPWR NMOS1_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0961_ _0413_ _0422_ VGND VPWR _0423_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_39_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0892_ _0370_ _0373_ VGND VPWR _0041_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_6_229 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1375_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0172_ VGND VPWR Dead_Time_Generator_inst_3.count_dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1091_ _0515_ VGND VPWR _0086_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1160_ _0208_ _0021_ _0211_ VGND VPWR _0537_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_67 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0944_ Shift_Register_Inst.data_out\[16\] net8 VGND VPWR _0411_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0875_ _0347_ _0359_ VGND VPWR _0360_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_2_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1358_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0045_ _0131_ VGND VPWR Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1289_ clknet_1_1__leaf_CLK_SR _0142_ _0063_ VGND VPWR Shift_Register_Inst.data_out\[10\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0660_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ Shift_Register_Inst.shift_state\[1\] VGND VPWR _0200_ VGND VPWR sky130_fd_sc_hd__or3b_2
X_1212_ Dead_Time_Generator_inst_2.count_dt\[0\] VGND VPWR _0583_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_46_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1143_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] VGND VPWR
+ _0520_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1074_ _0484_ _0491_ VGND VPWR _0508_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0927_ Signal_Generator_2_270phase_inst.count\[2\] _0392_ VGND VPWR _0399_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0858_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ VGND VPWR _0347_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0789_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR _0295_ VGND VPWR sky130_fd_sc_hd__o31ai_1
Xhold26 Signal_Generator_2_180phase_inst.direction VGND VPWR net51 VGND VPWR sky130_fd_sc_hd__buf_1
Xhold15 Dead_Time_Generator_inst_1.count_dt\[3\] VGND VPWR net40 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 Dead_Time_Generator_inst_3.count_dt\[2\] VGND VPWR net62 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0712_ _0183_ VGND VPWR _0237_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0643_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[1\]
+ Shift_Register_Inst.shift_state\[0\] VGND VPWR _0188_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1126_ _0518_ VGND VPWR _0118_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1057_ _0485_ _0489_ _0490_ VGND VPWR _0491_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_7_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput16 net16 VGND VPWR NMOS1_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1109_ _0516_ VGND VPWR _0103_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_23_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0960_ _0421_ net6 _0228_ VGND VPWR _0422_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0891_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0372_ VGND VPWR _0373_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_40_68 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1374_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0171_ VGND VPWR Dead_Time_Generator_inst_3.count_dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_122 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1090_ _0446_ VGND VPWR _0515_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_35_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0874_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VPWR _0359_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0943_ _0410_ VGND VPWR Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_0_2_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1288_ clknet_1_1__leaf_CLK_SR _0141_ _0062_ VGND VPWR Shift_Register_Inst.data_out\[11\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1357_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0044_ _0130_ VGND VPWR Signal_Generator_2_270phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1211_ Dead_Time_Generator_inst_2.count_dt\[1\] VGND VPWR _0582_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1142_ Shift_Register_Inst.data_out\[16\] net8 VGND VPWR _0519_ VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_46_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1073_ _0495_ _0496_ _0505_ _0506_ VGND VPWR _0507_ VGND VPWR sky130_fd_sc_hd__a211o_1
X_0926_ Signal_Generator_2_270phase_inst.count\[2\] _0395_ VGND VPWR _0398_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0857_ net65 Signal_Generator_2_0phase_inst.direction _0330_ _0346_ VGND VPWR _0033_
+ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_15_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0788_ _0285_ _0292_ _0294_ net55 VGND VPWR _0009_ VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold27 Signal_Generator_2_90phase_inst.direction VGND VPWR net52 VGND VPWR sky130_fd_sc_hd__buf_1
Xhold16 _0580_ VGND VPWR net41 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 Dead_Time_Generator_inst_1.count_dt\[2\] VGND VPWR net63 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0711_ _0236_ VGND VPWR _0136_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0642_ _0186_ _0187_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ net48 VGND VPWR _0156_ VGND VPWR sky130_fd_sc_hd__a41o_1
Xclkbuf_3_1__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_1125_ _0518_ VGND VPWR _0117_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1056_ Signal_Generator_2_0phase_inst.count\[2\] _0467_ VGND VPWR _0490_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0909_ Signal_Generator_2_180phase_inst.count\[4\] _0372_ VGND VPWR _0386_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
Xoutput17 net17 VGND VPWR NMOS2_PS1 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1108_ _0516_ VGND VPWR _0102_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1039_ _0214_ _0216_ Signal_Generator_2_270phase_inst.count\[5\] VGND VPWR _0473_
+ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_16_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0890_ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ _0371_ VGND VPWR _0372_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1373_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk net38 VGND VPWR Dead_Time_Generator_inst_3.count_dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_156 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0942_ CLK_PLL CLK_EXT Shift_Register_Inst.data_out\[14\] VGND VPWR _0410_ VGND VPWR
+ sky130_fd_sc_hd__mux2_4
X_0873_ _0349_ _0356_ _0358_ net52 VGND VPWR _0051_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_2_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1356_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0043_ _0129_ VGND VPWR Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1287_ clknet_1_1__leaf_CLK_SR _0140_ _0061_ VGND VPWR Shift_Register_Inst.data_out\[12\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1210_ _0447_ VGND VPWR _0134_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1141_ _0447_ VGND VPWR _0133_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1072_ _0502_ _0497_ _0501_ VGND VPWR _0506_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_46_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0856_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0326_ Signal_Generator_2_0phase_inst.count\[5\] VGND VPWR _0346_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0925_ _0048_ _0396_ _0397_ VGND VPWR _0043_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0787_ _0288_ _0293_ VGND VPWR _0294_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_30_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold17 Signal_Generator_1_0phase_inst.count\[0\] VGND VPWR net42 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 Signal_Generator_1_90phase_inst.count\[5\] VGND VPWR net53 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 Shift_Register_Inst.data_out\[15\] VGND VPWR net64 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1339_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0033_ _0112_ VGND VPWR Signal_Generator_2_0phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_0710_ net1 Shift_Register_Inst.data_out\[16\] _0235_ VGND VPWR _0236_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0641_ Shift_Register_Inst.shift_state\[2\] VGND VPWR _0187_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_1055_ _0471_ _0486_ _0487_ _0488_ VGND VPWR _0489_ VGND VPWR sky130_fd_sc_hd__or4_1
X_1124_ _0518_ VGND VPWR _0116_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0908_ _0382_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ VGND VPWR _0385_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0839_ _0332_ _0329_ VGND VPWR _0333_ VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput18 net18 VGND VPWR NMOS2_PS2 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1038_ Signal_Generator_2_90phase_inst.count\[5\] _0463_ _0464_ Signal_Generator_2_180phase_inst.count\[5\]
+ _0471_ VGND VPWR _0472_ VGND VPWR sky130_fd_sc_hd__a221o_1
X_1107_ _0516_ VGND VPWR _0101_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_17_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1372_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0169_ VGND VPWR Dead_Time_Generator_inst_1.go
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0941_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0393_ _0409_ VGND VPWR _0047_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0872_ _0352_ _0357_ VGND VPWR _0358_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1355_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0042_ _0128_ VGND VPWR Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1286_ clknet_1_0__leaf_CLK_SR _0139_ _0060_ VGND VPWR Shift_Register_Inst.data_out\[13\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1140_ _0447_ VGND VPWR _0132_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1071_ _0503_ _0504_ VGND VPWR _0505_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_46_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0924_ _0391_ _0396_ Signal_Generator_2_270phase_inst.direction VGND VPWR _0397_
+ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0786_ Signal_Generator_1_180phase_inst.count\[2\] _0286_ VGND VPWR _0293_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0855_ Signal_Generator_2_0phase_inst.direction _0343_ _0344_ _0328_ _0345_ VGND
+ VPWR _0032_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_30_108 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold18 Signal_Generator_1_90phase_inst.count\[0\] VGND VPWR net43 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 Signal_Generator_1_90phase_inst.direction VGND VPWR net54 VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
X_1338_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0032_ _0111_ VGND VPWR Signal_Generator_2_0phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1269_ Dead_Time_Generator_inst_4.count_dt\[1\] _0623_ VGND VPWR _0627_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_21_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_160 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_49 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0640_ Shift_Register_Inst.shift_state\[3\] VGND VPWR _0186_ VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_20_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1123_ _0446_ VGND VPWR _0518_ VGND VPWR sky130_fd_sc_hd__buf_4
X_1054_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_270phase_inst.count\[2\]
+ VGND VPWR _0488_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0907_ _0370_ _0381_ _0384_ net51 VGND VPWR _0038_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_7_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0769_ Signal_Generator_1_90phase_inst.count\[4\] _0261_ VGND VPWR _0281_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0838_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VPWR _0332_ VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput19 net19 VGND VPWR NMOS_PS3 VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1106_ _0516_ VGND VPWR _0100_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1037_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] VGND VPWR
+ _0471_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_17_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1371_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0168_ VGND VPWR Dead_Time_Generator_inst_2.count_dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0940_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0389_ Signal_Generator_2_270phase_inst.count\[5\] VGND VPWR _0409_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0871_ Signal_Generator_2_90phase_inst.count\[2\] _0350_ VGND VPWR _0357_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1285_ clknet_1_0__leaf_CLK_SR _0138_ _0059_ VGND VPWR Shift_Register_Inst.data_out\[14\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1354_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0048_ _0127_ VGND VPWR Signal_Generator_2_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1070_ _0495_ _0496_ VGND VPWR _0504_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0854_ Signal_Generator_2_0phase_inst.count\[4\] _0326_ VGND VPWR _0345_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0923_ _0395_ _0392_ VGND VPWR _0396_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_11_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0785_ Signal_Generator_1_180phase_inst.count\[2\] _0289_ VGND VPWR _0292_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_150 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1268_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_4.count_dt\[0\]
+ _0461_ VGND VPWR _0626_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1337_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0031_ _0110_ VGND VPWR Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xhold19 Signal_Generator_1_180phase_inst.count\[0\] VGND VPWR net44 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1199_ _0561_ _0574_ _0575_ VGND VPWR _0158_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_14_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1122_ _0517_ VGND VPWR _0115_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1053_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[2\]
+ Shift_Register_Inst.data_out\[7\] VGND VPWR _0487_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0906_ _0382_ _0383_ _0373_ VGND VPWR _0384_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0837_ net34 VGND VPWR _0028_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_94 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0768_ Signal_Generator_1_90phase_inst.count\[4\] _0266_ VGND VPWR _0280_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0699_ Shift_Register_Inst.data_out\[13\] VGND VPWR _0228_ VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_34_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1105_ _0516_ VGND VPWR _0099_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1036_ net14 VGND VPWR _0470_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_31_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1019_ Dead_Time_Generator_inst_4.count_dt\[0\] VGND VPWR _0453_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1370_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0167_ VGND VPWR Dead_Time_Generator_inst_2.count_dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0870_ Signal_Generator_2_90phase_inst.count\[2\] _0353_ VGND VPWR _0356_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
Xclkbuf_3_2__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_1284_ clknet_1_0__leaf_CLK_SR _0137_ _0058_ VGND VPWR Shift_Register_Inst.data_out\[15\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1353_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0040_ _0126_ VGND VPWR Signal_Generator_2_180phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_0999_ _0448_ VGND VPWR _0062_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_33_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0853_ Signal_Generator_2_0phase_inst.count\[4\] _0330_ VGND VPWR _0344_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0922_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VPWR _0395_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0784_ _0013_ _0290_ _0291_ VGND VPWR _0008_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1198_ net56 _0573_ VGND VPWR _0575_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1267_ _0625_ VGND VPWR _0176_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput1 Data_SR VGND VPWR net1 VGND VPWR sky130_fd_sc_hd__buf_2
X_1336_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0030_ _0109_ VGND VPWR Signal_Generator_2_0phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1121_ _0517_ VGND VPWR _0114_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1052_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_180phase_inst.count\[2\]
+ VGND VPWR _0486_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_7_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0767_ _0276_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ VGND VPWR _0279_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0905_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VPWR _0383_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0836_ _0328_ _0331_ VGND VPWR _0034_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0698_ _0227_ VGND VPWR _0140_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1319_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0013_ _0092_ VGND VPWR Signal_Generator_1_180phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1104_ _0516_ VGND VPWR _0098_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1035_ _0462_ _0468_ VGND VPWR _0469_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_17_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0819_ _0305_ _0317_ VGND VPWR _0318_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_31_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1018_ Dead_Time_Generator_inst_4.count_dt\[1\] VGND VPWR _0452_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1352_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0039_ _0125_ VGND VPWR Signal_Generator_2_180phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1283_ clknet_1_0__leaf_CLK_SR _0136_ _0057_ VGND VPWR Shift_Register_Inst.data_out\[16\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0998_ _0448_ VGND VPWR _0061_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_33_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0921_ net32 VGND VPWR _0042_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0852_ _0340_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ VGND VPWR _0343_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0783_ _0285_ _0290_ net55 VGND VPWR _0291_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_86 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1335_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0029_ _0108_ VGND VPWR Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1197_ Dead_Time_Generator_inst_1.count_dt\[0\] _0573_ VGND VPWR _0574_ VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1266_ _0623_ _0624_ _0513_ VGND VPWR _0625_ VGND VPWR sky130_fd_sc_hd__and3b_1
Xinput2 RST VGND VPWR net2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_166 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1120_ _0517_ VGND VPWR _0113_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1051_ net11 VGND VPWR _0485_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0904_ _0372_ VGND VPWR _0382_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_22_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0697_ net1 Shift_Register_Inst.data_out\[12\] _0226_ VGND VPWR _0227_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0766_ _0263_ _0275_ _0278_ net54 VGND VPWR _0024_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0835_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0330_ VGND VPWR _0331_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1318_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0026_ _0091_ VGND VPWR Signal_Generator_1_90phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1249_ net27 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VPWR _0614_ VGND VPWR
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1034_ Signal_Generator_2_0phase_inst.count\[4\] _0466_ _0467_ VGND VPWR _0468_ VGND
+ VPWR sky130_fd_sc_hd__mux2_1
X_1103_ _0516_ VGND VPWR _0097_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_31_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0818_ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR _0317_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0749_ _0264_ _0021_ VGND VPWR _0265_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_38_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1017_ Dead_Time_Generator_inst_4.count_dt\[2\] VGND VPWR _0451_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1351_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0038_ _0124_ VGND VPWR Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1282_ clknet_1_0__leaf_CLK_SR _0135_ _0056_ VGND VPWR Shift_Register_Inst.data_out\[17\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0997_ _0448_ VGND VPWR _0060_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_41_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0920_ _0391_ _0394_ VGND VPWR _0048_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0851_ _0328_ _0339_ _0342_ Signal_Generator_2_0phase_inst.direction VGND VPWR _0031_
+ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0782_ _0289_ _0286_ VGND VPWR _0290_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_11_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1265_ Dead_Time_Generator_inst_4.count_dt\[0\] _0461_ VGND VPWR _0624_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1334_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0028_ _0107_ VGND VPWR Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1196_ _0569_ _0570_ _0571_ _0572_ VGND VPWR _0573_ VGND VPWR sky130_fd_sc_hd__o31a_1
Xinput3 d1[0] VGND VPWR net3 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_14_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1050_ _0478_ _0482_ _0483_ VGND VPWR _0484_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0903_ _0368_ _0380_ VGND VPWR _0381_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0834_ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ _0329_ VGND VPWR _0330_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_43_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0765_ _0276_ _0277_ _0267_ VGND VPWR _0278_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0696_ _0225_ _0205_ VGND VPWR _0226_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1248_ Dead_Time_Generator_inst_3.count_dt\[4\] net27 VGND VPWR _0613_ VGND VPWR
+ sky130_fd_sc_hd__and2b_1
X_1317_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0025_ _0090_ VGND VPWR Signal_Generator_1_90phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1179_ _0551_ _0552_ VGND VPWR _0556_ VGND VPWR sky130_fd_sc_hd__nand2_1
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1102_ _0516_ VGND VPWR _0096_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1033_ _0214_ _0216_ VGND VPWR _0467_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0817_ _0307_ _0314_ _0316_ Signal_Generator_1_270phase_inst.direction VGND VPWR
+ _0016_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_24_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0748_ net43 VGND VPWR _0021_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0679_ Shift_Register_Inst.data_out\[7\] VGND VPWR _0214_ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1016_ _0450_ VGND VPWR _0077_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_8_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1281_ _0513_ net29 VGND VPWR _0181_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1350_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0037_ _0123_ VGND VPWR Signal_Generator_2_180phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_0996_ _0448_ VGND VPWR _0059_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_1_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0850_ _0340_ _0341_ _0331_ VGND VPWR _0342_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0781_ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VPWR _0289_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1264_ Dead_Time_Generator_inst_4.count_dt\[0\] _0461_ VGND VPWR _0623_ VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1333_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0034_ _0106_ VGND VPWR Signal_Generator_2_0phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
Xinput4 d1[1] VGND VPWR net4 VGND VPWR sky130_fd_sc_hd__buf_1
X_1195_ net27 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VPWR _0572_ VGND VPWR
+ sky130_fd_sc_hd__or2b_1
X_0979_ net20 _0430_ _0433_ _0435_ Shift_Register_Inst.data_out\[11\] VGND VPWR _0436_
+ VGND VPWR sky130_fd_sc_hd__a2111o_1
X_0902_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VPWR _0380_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0833_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ VGND VPWR _0329_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_43_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0695_ _0186_ _0187_ VGND VPWR _0225_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0764_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VPWR _0277_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_11_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1178_ _0535_ _0541_ _0554_ VGND VPWR _0555_ VGND VPWR sky130_fd_sc_hd__o21ai_1
X_1247_ _0609_ Dead_Time_Generator_inst_1.dt\[3\] VGND VPWR _0612_ VGND VPWR sky130_fd_sc_hd__and2_1
X_1316_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0024_ _0089_ VGND VPWR Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1032_ Signal_Generator_2_90phase_inst.count\[4\] _0463_ _0464_ Signal_Generator_2_180phase_inst.count\[4\]
+ _0465_ VGND VPWR _0466_ VGND VPWR sky130_fd_sc_hd__a221o_1
X_1101_ _0446_ VGND VPWR _0516_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_33_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0747_ Signal_Generator_1_90phase_inst.count\[1\] VGND VPWR _0264_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0816_ _0310_ _0315_ VGND VPWR _0316_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_16_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0678_ _0213_ VGND VPWR _0146_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1015_ _0450_ VGND VPWR _0076_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_30_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1280_ net30 _0632_ _0513_ VGND VPWR _0180_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_25_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0995_ _0448_ VGND VPWR _0058_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0780_ net44 VGND VPWR _0007_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1194_ Dead_Time_Generator_inst_1.count_dt\[4\] net27 VGND VPWR _0571_ VGND VPWR
+ sky130_fd_sc_hd__and2b_1
X_1263_ _0581_ _0593_ VGND VPWR _0175_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1332_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0019_ _0105_ VGND VPWR Signal_Generator_1_270phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
Xinput5 d1[2] VGND VPWR net5 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_46_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0978_ _0431_ net15 _0434_ Shift_Register_Inst.data_out\[10\] VGND VPWR _0435_ VGND
+ VPWR sky130_fd_sc_hd__o211a_1
X_0901_ _0370_ _0377_ _0379_ net51 VGND VPWR _0037_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0763_ _0266_ VGND VPWR _0276_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0832_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0326_ _0327_ VGND VPWR _0328_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_1315_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0023_ _0088_ VGND VPWR Signal_Generator_1_90phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_0_11_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0694_ _0224_ VGND VPWR _0141_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1177_ _0551_ _0552_ _0553_ VGND VPWR _0554_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1246_ _0606_ _0608_ _0610_ VGND VPWR _0611_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_33_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1100_ _0515_ VGND VPWR _0095_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1031_ _0214_ _0216_ Signal_Generator_2_270phase_inst.count\[4\] VGND VPWR _0465_
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_0746_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0261_ _0262_ VGND VPWR _0263_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_0815_ Signal_Generator_1_270phase_inst.count\[2\] _0308_ VGND VPWR _0315_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0677_ _0182_ _0211_ _0212_ VGND VPWR _0213_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1229_ _0597_ _0598_ _0561_ VGND VPWR _0599_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_30_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1014_ _0446_ VGND VPWR _0450_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_44_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0729_ Signal_Generator_1_0phase_inst.count\[2\] _0243_ VGND VPWR _0250_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0994_ _0448_ VGND VPWR _0057_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1331_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0018_ _0104_ VGND VPWR Signal_Generator_1_270phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1262_ net33 _0621_ _0513_ VGND VPWR _0174_ VGND VPWR sky130_fd_sc_hd__o21ba_1
X_1193_ _0567_ net39 VGND VPWR _0570_ VGND VPWR sky130_fd_sc_hd__and2_1
Xinput6 d1[3] VGND VPWR net6 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_46_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0977_ Shift_Register_Inst.data_out\[9\] net22 VGND VPWR _0434_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_9_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0900_ _0373_ _0378_ VGND VPWR _0379_ VGND VPWR sky130_fd_sc_hd__or2_1
XPHY_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0693_ Shift_Register_Inst.data_out\[11\] net1 _0223_ VGND VPWR _0224_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0831_ Signal_Generator_2_0phase_inst.direction VGND VPWR _0327_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0762_ _0261_ _0274_ VGND VPWR _0275_ VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_0_11_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_Dead_Time_Generator_inst_1.clk Dead_Time_Generator_inst_1.clk VGND VPWR
+ clknet_0_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_1314_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0022_ _0087_ VGND VPWR Signal_Generator_1_90phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1245_ _0607_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0609_ VGND VPWR _0610_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1176_ _0549_ _0550_ VGND VPWR _0553_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_42_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1030_ _0214_ _0216_ VGND VPWR _0464_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0814_ Signal_Generator_1_270phase_inst.count\[2\] _0311_ VGND VPWR _0314_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0676_ _0200_ _0186_ Shift_Register_Inst.shift_state\[2\] VGND VPWR _0212_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_0745_ Signal_Generator_1_90phase_inst.direction VGND VPWR _0262_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1228_ Dead_Time_Generator_inst_2.count_dt\[1\] _0594_ VGND VPWR _0598_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1159_ _0208_ _0211_ Signal_Generator_1_270phase_inst.count\[0\] VGND VPWR _0536_
+ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_30_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1013_ _0449_ VGND VPWR _0075_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0728_ Signal_Generator_1_0phase_inst.count\[2\] _0246_ VGND VPWR _0249_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0659_ _0199_ VGND VPWR _0151_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_187 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0993_ _0448_ VGND VPWR _0056_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_1_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1261_ _0513_ _0621_ _0622_ VGND VPWR _0173_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1330_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0017_ _0103_ VGND VPWR Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1192_ _0564_ _0566_ _0568_ VGND VPWR _0569_ VGND VPWR sky130_fd_sc_hd__o21a_1
Xinput7 d1[4] VGND VPWR net7 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_36_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0976_ net17 _0432_ VGND VPWR _0433_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_46_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_190 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0830_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ VGND VPWR _0326_ VGND VPWR sky130_fd_sc_hd__or4_2
XPHY_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0761_ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VPWR _0274_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0692_ _0187_ _0188_ _0186_ VGND VPWR _0223_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1244_ Dead_Time_Generator_inst_3.count_dt\[3\] VGND VPWR _0609_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1313_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0021_ _0086_ VGND VPWR Signal_Generator_1_90phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1175_ _0547_ _0548_ _0542_ VGND VPWR _0552_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0959_ Dead_Time_Generator_inst_1.go VGND VPWR _0421_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_6_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0813_ _0020_ _0312_ _0313_ VGND VPWR _0015_ VGND VPWR sky130_fd_sc_hd__a21oi_1
Xinput10 d2[1] VGND VPWR net10 VGND VPWR sky130_fd_sc_hd__buf_1
X_0744_ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ Signal_Generator_1_90phase_inst.count\[1\] Signal_Generator_1_90phase_inst.count\[0\]
+ VGND VPWR _0261_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0675_ Shift_Register_Inst.data_out\[6\] VGND VPWR _0211_ VGND VPWR sky130_fd_sc_hd__buf_2
X_1227_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_2.count_dt\[0\]
+ _0593_ VGND VPWR _0597_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1158_ _0228_ _0530_ _0534_ VGND VPWR _0535_ VGND VPWR sky130_fd_sc_hd__o21a_1
X_1089_ _0450_ VGND VPWR _0085_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1012_ _0449_ VGND VPWR _0074_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0727_ _0006_ _0247_ _0248_ VGND VPWR _0001_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0658_ _0182_ Dead_Time_Generator_inst_1.dt\[1\] _0198_ VGND VPWR _0199_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_199 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0992_ _0447_ VGND VPWR _0448_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_41_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1191_ _0565_ Dead_Time_Generator_inst_1.dt\[2\] Dead_Time_Generator_inst_1.dt\[3\]
+ _0567_ VGND VPWR _0568_ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1260_ Dead_Time_Generator_inst_3.count_dt\[2\] _0618_ net45 VGND VPWR _0622_ VGND
+ VPWR sky130_fd_sc_hd__a21oi_1
Xinput8 d1[5] VGND VPWR net8 VGND VPWR sky130_fd_sc_hd__buf_1
X_0975_ _0431_ Shift_Register_Inst.data_out\[10\] VGND VPWR _0432_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_45_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_0760_ _0263_ _0271_ _0273_ net54 VGND VPWR _0023_ VGND VPWR sky130_fd_sc_hd__a22o_1
XPHY_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0691_ _0222_ VGND VPWR _0142_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1174_ _0542_ _0547_ _0548_ _0549_ _0550_ VGND VPWR _0551_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_1243_ _0604_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[2\]
+ _0607_ VGND VPWR _0608_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_1312_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0027_ _0085_ VGND VPWR Signal_Generator_1_90phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_19_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0889_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ VGND VPWR _0371_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0958_ _0420_ VGND VPWR net18 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_34_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_161 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0812_ _0307_ _0312_ Signal_Generator_1_270phase_inst.direction VGND VPWR _0313_
+ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0743_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0244_ _0260_ VGND VPWR _0005_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xinput11 d2[2] VGND VPWR net11 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0674_ _0210_ VGND VPWR _0147_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1157_ Signal_Generator_1_0phase_inst.count\[1\] _0520_ _0532_ _0533_ VGND VPWR _0534_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
X_1226_ _0596_ VGND VPWR _0164_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1088_ _0450_ VGND VPWR _0084_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_2_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1011_ _0449_ VGND VPWR _0073_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0726_ _0242_ _0247_ net58 VGND VPWR _0248_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0657_ Shift_Register_Inst.shift_state\[4\] _0194_ _0183_ VGND VPWR _0198_ VGND VPWR
+ sky130_fd_sc_hd__or3_1
XFILLER_0_33_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1209_ net36 _0579_ _0581_ VGND VPWR _0162_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_30_47 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0709_ Shift_Register_Inst.shift_state\[0\] _0183_ Shift_Register_Inst.shift_state\[4\]
+ VGND VPWR _0235_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_4_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0991_ _0446_ VGND VPWR _0447_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_41_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1190_ Dead_Time_Generator_inst_1.count_dt\[3\] VGND VPWR _0567_ VGND VPWR sky130_fd_sc_hd__inv_2
Xinput9 d2[0] VGND VPWR net9 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0974_ Shift_Register_Inst.data_out\[9\] VGND VPWR _0431_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_14_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0690_ net1 Shift_Register_Inst.data_out\[10\] _0221_ VGND VPWR _0222_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1311_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0005_ _0084_ VGND VPWR Signal_Generator_1_0phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1173_ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[2\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[2\]
+ Shift_Register_Inst.data_out\[5\] _0211_ VGND VPWR _0550_ VGND VPWR sky130_fd_sc_hd__mux4_1
X_1242_ Dead_Time_Generator_inst_3.count_dt\[2\] VGND VPWR _0607_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_27_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0413_ _0419_ VGND VPWR _0420_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0888_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0368_ _0369_ VGND VPWR _0370_ VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_42_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_173 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0673_ _0182_ _0208_ _0209_ VGND VPWR _0210_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0742_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0240_ Signal_Generator_1_0phase_inst.count\[5\] VGND VPWR _0260_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0811_ _0311_ _0308_ VGND VPWR _0312_ VGND VPWR sky130_fd_sc_hd__or2_1
Xinput12 d2[3] VGND VPWR net12 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1087_ _0450_ VGND VPWR _0083_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1156_ _0208_ _0264_ _0211_ VGND VPWR _0533_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1225_ _0594_ _0595_ _0561_ VGND VPWR _0596_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_28_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1010_ _0449_ VGND VPWR _0072_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0656_ net60 _0195_ VGND VPWR _0152_ VGND VPWR sky130_fd_sc_hd__xnor2_1
X_0725_ _0246_ _0243_ VGND VPWR _0247_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_8_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1208_ _0529_ _0558_ _0559_ _0560_ VGND VPWR _0581_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_26_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1139_ _0447_ VGND VPWR _0131_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0639_ _0185_ VGND VPWR _0163_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0708_ _0234_ VGND VPWR _0137_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0990_ net2 VGND VPWR _0446_ VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0973_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] VGND
+ VPWR _0430_ VGND VPWR sky130_fd_sc_hd__nor2_1
XPHY_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1241_ _0604_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[0\]
+ _0605_ VGND VPWR _0606_ VGND VPWR sky130_fd_sc_hd__o211a_1
X_1310_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0004_ _0083_ VGND VPWR Signal_Generator_1_0phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1172_ _0228_ net5 VGND VPWR _0549_ VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0956_ Dead_Time_Generator_inst_2.go net3 _0228_ VGND VPWR _0419_ VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_27_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0887_ Signal_Generator_2_180phase_inst.direction VGND VPWR _0369_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_33_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0810_ Signal_Generator_1_270phase_inst.count\[1\] Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR _0311_ VGND VPWR sky130_fd_sc_hd__nor2_1
Xinput13 d2[4] VGND VPWR net13 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0672_ _0196_ _0186_ Shift_Register_Inst.shift_state\[2\] VGND VPWR _0209_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_0741_ Signal_Generator_1_0phase_inst.direction _0257_ _0258_ _0242_ _0259_ VGND
+ VPWR _0004_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_1224_ Dead_Time_Generator_inst_2.count_dt\[0\] _0593_ VGND VPWR _0595_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1086_ _0450_ VGND VPWR _0082_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1155_ _0208_ _0211_ Signal_Generator_1_270phase_inst.count\[1\] _0531_ VGND VPWR
+ _0532_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0939_ Signal_Generator_2_270phase_inst.direction _0406_ _0407_ _0391_ _0408_ VGND
+ VPWR _0046_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_23_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0655_ _0196_ _0197_ VGND VPWR _0153_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0724_ Signal_Generator_1_0phase_inst.count\[1\] Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VPWR _0246_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_12_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1207_ _0561_ _0579_ net41 VGND VPWR _0161_ VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_0_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1069_ _0497_ _0501_ _0502_ VGND VPWR _0503_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_1138_ _0447_ VGND VPWR _0130_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_252 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold2 Dead_Time_Generator_inst_1.dt\[4\] VGND VPWR net27 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_0707_ net64 net1 _0233_ VGND VPWR _0234_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_0638_ _0182_ Dead_Time_Generator_inst_1.dt\[0\] _0184_ VGND VPWR _0185_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0972_ Shift_Register_Inst.data_out\[12\] VGND VPWR _0429_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_39_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1240_ Dead_Time_Generator_inst_3.count_dt\[0\] VGND VPWR _0605_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1171_ Signal_Generator_1_0phase_inst.count\[3\] _0520_ VGND VPWR _0548_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0886_ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ VGND VPWR _0368_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0955_ _0418_ VGND VPWR net23 VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_1369_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0166_ VGND VPWR Dead_Time_Generator_inst_2.count_dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0740_ Signal_Generator_1_0phase_inst.count\[4\] _0240_ VGND VPWR _0259_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
Xinput14 d2[5] VGND VPWR net14 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0671_ Shift_Register_Inst.data_out\[5\] VGND VPWR _0208_ VGND VPWR sky130_fd_sc_hd__buf_2
X_1223_ Dead_Time_Generator_inst_2.count_dt\[0\] _0593_ VGND VPWR _0594_ VGND VPWR
+ sky130_fd_sc_hd__and2_1
X_1154_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VPWR _0531_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1085_ _0450_ VGND VPWR _0081_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0938_ Signal_Generator_2_270phase_inst.count\[4\] _0389_ VGND VPWR _0408_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0869_ _0055_ _0354_ _0355_ VGND VPWR _0050_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0723_ net42 VGND VPWR _0000_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0654_ net48 _0194_ net57 VGND VPWR _0197_ VGND VPWR sky130_fd_sc_hd__o21ai_1
X_1137_ _0447_ VGND VPWR _0129_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1206_ Dead_Time_Generator_inst_1.count_dt\[2\] _0576_ net40 VGND VPWR _0580_ VGND
+ VPWR sky130_fd_sc_hd__a21oi_1
X_1068_ net10 VGND VPWR _0502_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold3 _0614_ VGND VPWR net28 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0706_ _0186_ _0187_ _0188_ VGND VPWR _0233_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0637_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ _0183_ VGND VPWR _0184_ VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_0_29_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_5__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0971_ _0428_ VGND VPWR net20 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_39_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1170_ _0543_ _0544_ _0545_ _0546_ VGND VPWR _0547_ VGND VPWR sky130_fd_sc_hd__or4_1
X_0954_ _0413_ _0416_ _0417_ VGND VPWR _0418_ VGND VPWR sky130_fd_sc_hd__or3_1
X_0885_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0351_ _0367_ VGND VPWR _0054_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_1368_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0165_ VGND VPWR Dead_Time_Generator_inst_2.count_dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1299_ clknet_1_0__leaf_CLK_SR _0152_ _0073_ VGND VPWR Shift_Register_Inst.shift_state\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0670_ _0207_ VGND VPWR _0148_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1153_ net4 VGND VPWR _0530_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1084_ _0450_ VGND VPWR _0080_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1222_ _0589_ _0590_ _0591_ _0592_ VGND VPWR _0593_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0799_ _0301_ _0302_ _0285_ _0303_ VGND VPWR _0011_ VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_0868_ _0349_ _0354_ net52 VGND VPWR _0355_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0937_ Signal_Generator_2_270phase_inst.count\[4\] _0393_ VGND VPWR _0407_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0653_ Shift_Register_Inst.shift_state\[1\] _0194_ _0195_ VGND VPWR _0196_ VGND VPWR
+ sky130_fd_sc_hd__or3_2
X_0722_ _0242_ _0245_ VGND VPWR _0006_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1067_ _0471_ _0498_ _0499_ _0500_ VGND VPWR _0501_ VGND VPWR sky130_fd_sc_hd__or4_1
X_1136_ _0447_ VGND VPWR _0128_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1205_ Dead_Time_Generator_inst_1.count_dt\[3\] Dead_Time_Generator_inst_1.count_dt\[2\]
+ _0576_ VGND VPWR _0579_ VGND VPWR sky130_fd_sc_hd__and3_1
Xhold4 _0615_ VGND VPWR net29 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0636_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ Shift_Register_Inst.shift_state\[1\] VGND VPWR _0183_ VGND VPWR sky130_fd_sc_hd__or3_2
X_0705_ _0232_ VGND VPWR _0138_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1119_ _0517_ VGND VPWR _0112_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_0_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_17 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0970_ _0422_ _0424_ VGND VPWR _0428_ VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_26_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1384_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0181_ VGND VPWR Dead_Time_Generator_inst_3.go
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_60 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0884_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0347_ Signal_Generator_2_90phase_inst.count\[5\] VGND VPWR _0367_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0953_ _0228_ Dead_Time_Generator_inst_3.go VGND VPWR _0417_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_12_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1367_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0164_ VGND VPWR Dead_Time_Generator_inst_2.count_dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1298_ clknet_1_0__leaf_CLK_SR _0151_ _0072_ VGND VPWR Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1221_ net27 Dead_Time_Generator_inst_2.count_dt\[4\] VGND VPWR _0592_ VGND VPWR
+ sky130_fd_sc_hd__or2b_1
Xclkbuf_1_1__f_CLK_SR clknet_0_CLK_SR VGND VPWR clknet_1_1__leaf_CLK_SR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_1083_ _0450_ VGND VPWR _0079_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1152_ _0525_ _0528_ VGND VPWR _0529_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0936_ _0403_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VPWR _0406_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_15_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0798_ Signal_Generator_1_180phase_inst.count\[4\] _0283_ VGND VPWR _0303_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0867_ _0353_ _0350_ VGND VPWR _0354_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_15_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0652_ Shift_Register_Inst.shift_state\[4\] _0183_ VGND VPWR _0195_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0721_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0244_ VGND VPWR _0245_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1204_ _0561_ _0578_ VGND VPWR _0160_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_20_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1135_ _0447_ VGND VPWR _0127_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1066_ _0214_ _0216_ Signal_Generator_2_270phase_inst.count\[1\] VGND VPWR _0500_
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_0919_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0393_ VGND VPWR _0394_ VGND VPWR sky130_fd_sc_hd__and3_1
Xhold5 Dead_Time_Generator_inst_4.count_dt\[4\] VGND VPWR net30 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0704_ net1 Shift_Register_Inst.data_out\[14\] _0231_ VGND VPWR _0232_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0635_ net1 VGND VPWR _0182_ VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_17_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_71 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1118_ _0517_ VGND VPWR _0111_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1049_ Signal_Generator_2_0phase_inst.count\[3\] _0467_ VGND VPWR _0483_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_34_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1383_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0180_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0952_ _0228_ net4 VGND VPWR _0416_ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_42_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0883_ net52 _0364_ _0365_ _0349_ _0366_ VGND VPWR _0053_ VGND VPWR sky130_fd_sc_hd__a32o_1
XFILLER_0_12_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1366_ clknet_1_0__leaf_CLK_SR _0163_ _0134_ VGND VPWR Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1297_ clknet_1_0__leaf_CLK_SR _0150_ _0071_ VGND VPWR Dead_Time_Generator_inst_1.dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1151_ _0519_ _0524_ _0526_ _0527_ VGND VPWR _0528_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_1220_ Dead_Time_Generator_inst_2.count_dt\[4\] net27 VGND VPWR _0591_ VGND VPWR
+ sky130_fd_sc_hd__and2b_1
X_1082_ _0450_ VGND VPWR _0078_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0935_ _0391_ _0402_ _0405_ Signal_Generator_2_270phase_inst.direction VGND VPWR
+ _0045_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0866_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ VGND VPWR _0353_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_15_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0797_ Signal_Generator_1_180phase_inst.count\[4\] _0287_ Signal_Generator_1_180phase_inst.direction
+ VGND VPWR _0302_ VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1349_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0036_ _0122_ VGND VPWR Signal_Generator_2_180phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0720_ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ _0243_ VGND VPWR _0244_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0651_ Shift_Register_Inst.shift_state\[0\] VGND VPWR _0194_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1134_ _0447_ VGND VPWR _0126_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1203_ net63 _0576_ VGND VPWR _0578_ VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_52 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1065_ _0214_ _0216_ Signal_Generator_2_180phase_inst.count\[1\] VGND VPWR _0499_
+ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0918_ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ _0392_ VGND VPWR _0393_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0849_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR _0341_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_11_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold6 Dead_Time_Generator_inst_2.count_dt\[4\] VGND VPWR net31 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0703_ _0225_ _0200_ VGND VPWR _0231_ VGND VPWR sky130_fd_sc_hd__or2_1
X_1117_ _0517_ VGND VPWR _0110_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_45_83 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1048_ _0471_ _0479_ _0480_ _0481_ VGND VPWR _0482_ VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_0_28_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_63 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1382_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0179_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0882_ Signal_Generator_2_90phase_inst.count\[4\] _0347_ VGND VPWR _0366_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0951_ _0415_ VGND VPWR net16 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_42_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1365_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0162_ VGND VPWR Dead_Time_Generator_inst_1.count_dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1296_ clknet_1_0__leaf_CLK_SR _0149_ _0070_ VGND VPWR Dead_Time_Generator_inst_1.dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1150_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_90phase_inst.count\[4\]
+ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0208_ _0211_ VGND VPWR _0527_ VGND VPWR sky130_fd_sc_hd__mux4_1
X_1081_ _0514_ VGND VPWR _0157_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0934_ _0403_ _0404_ _0394_ VGND VPWR _0405_ VGND VPWR sky130_fd_sc_hd__a21o_1
X_0865_ net46 VGND VPWR _0049_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_15_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6__f_Dead_Time_Generator_inst_1.clk net26 VGND VPWR clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_0796_ _0300_ Signal_Generator_1_180phase_inst.count\[4\] _0287_ VGND VPWR _0301_
+ VGND VPWR sky130_fd_sc_hd__and3_1
X_1348_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0035_ _0121_ VGND VPWR Signal_Generator_2_180phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1279_ _0634_ VGND VPWR _0179_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0650_ _0193_ VGND VPWR _0154_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1133_ _0518_ VGND VPWR _0125_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1202_ _0561_ _0576_ _0577_ VGND VPWR _0159_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1064_ _0216_ Signal_Generator_2_90phase_inst.count\[1\] _0214_ VGND VPWR _0498_
+ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_18_64 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0848_ _0330_ VGND VPWR _0340_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0917_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ VGND VPWR _0392_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0779_ _0285_ _0288_ VGND VPWR _0013_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_11_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_CLK_SR CLK_SR VGND VPWR clknet_0_CLK_SR VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold7 Signal_Generator_2_270phase_inst.count\[0\] VGND VPWR net32 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0702_ _0230_ VGND VPWR _0139_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1116_ _0517_ VGND VPWR _0109_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1047_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR _0481_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_45_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1381_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0178_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_149 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0950_ _0413_ _0414_ VGND VPWR _0415_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0881_ Signal_Generator_2_90phase_inst.count\[4\] _0351_ VGND VPWR _0365_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_12_55 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1295_ clknet_1_0__leaf_CLK_SR _0148_ _0069_ VGND VPWR Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1364_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0161_ VGND VPWR Dead_Time_Generator_inst_1.count_dt\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1080_ _0461_ _0513_ VGND VPWR _0514_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0795_ Signal_Generator_1_180phase_inst.count\[5\] VGND VPWR _0300_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0933_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR _0404_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0864_ _0349_ _0352_ VGND VPWR _0055_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1347_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0041_ _0120_ VGND VPWR Signal_Generator_2_180phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1278_ _0632_ _0633_ _0512_ VGND VPWR _0634_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1201_ net49 _0574_ VGND VPWR _0577_ VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_0_20_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1132_ _0518_ VGND VPWR _0124_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1063_ Signal_Generator_2_0phase_inst.count\[1\] _0467_ VGND VPWR _0497_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_0916_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0389_ _0390_ VGND VPWR _0391_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0847_ _0326_ _0338_ VGND VPWR _0339_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0778_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0287_ VGND VPWR _0288_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_11_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold8 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VPWR net33 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0701_ net1 _0228_ _0229_ VGND VPWR _0230_ VGND VPWR sky130_fd_sc_hd__mux2_1
X_1115_ _0517_ VGND VPWR _0108_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1046_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[3\]
+ Shift_Register_Inst.data_out\[7\] VGND VPWR _0480_ VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_0_3_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1029_ _0216_ _0214_ VGND VPWR _0463_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_1380_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0177_ VGND VPWR Dead_Time_Generator_inst_4.count_dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0880_ _0361_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ VGND VPWR _0364_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_6_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1363_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0160_ VGND VPWR Dead_Time_Generator_inst_1.count_dt\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_1294_ clknet_1_1__leaf_CLK_SR _0147_ _0068_ VGND VPWR Shift_Register_Inst.data_out\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0932_ _0393_ VGND VPWR _0403_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0794_ _0285_ _0296_ _0299_ net55 VGND VPWR _0010_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0863_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0351_ VGND VPWR _0352_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1346_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0054_ _0119_ VGND VPWR Signal_Generator_2_90phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_1277_ Dead_Time_Generator_inst_4.count_dt\[2\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ _0623_ Dead_Time_Generator_inst_4.count_dt\[3\] VGND VPWR _0633_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_14_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1200_ Dead_Time_Generator_inst_1.count_dt\[1\] Dead_Time_Generator_inst_1.count_dt\[0\]
+ _0573_ VGND VPWR _0576_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1062_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[0\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[0\]
+ _0214_ _0216_ VGND VPWR _0496_ VGND VPWR sky130_fd_sc_hd__mux4_1
X_1131_ _0518_ VGND VPWR _0123_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_34_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0915_ Signal_Generator_2_270phase_inst.direction VGND VPWR _0390_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0846_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VPWR _0338_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0777_ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ _0286_ VGND VPWR _0287_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_45_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1329_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0016_ _0102_ VGND VPWR Signal_Generator_1_270phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold9 Signal_Generator_2_0phase_inst.count\[0\] VGND VPWR net34 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ _0225_ _0196_ VGND VPWR _0229_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_4_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1114_ _0517_ VGND VPWR _0107_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_45_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1045_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VPWR _0479_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_0829_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0309_ _0325_ VGND VPWR _0019_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_9_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1028_ net13 VGND VPWR _0462_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_16_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1293_ clknet_1_1__leaf_CLK_SR _0146_ _0067_ VGND VPWR Shift_Register_Inst.data_out\[6\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1362_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0159_ VGND VPWR Dead_Time_Generator_inst_1.count_dt\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0931_ _0389_ _0401_ VGND VPWR _0402_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_0862_ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ _0350_ VGND VPWR _0351_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0793_ _0297_ _0298_ _0288_ VGND VPWR _0299_ VGND VPWR sky130_fd_sc_hd__a21o_1
Xrebuffer1 clknet_0_Dead_Time_Generator_inst_1.clk VGND VPWR net26 VGND VPWR sky130_fd_sc_hd__buf_8
X_1276_ Dead_Time_Generator_inst_4.count_dt\[3\] Dead_Time_Generator_inst_4.count_dt\[2\]
+ _0626_ VGND VPWR _0632_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1345_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0053_ _0118_ VGND VPWR Signal_Generator_2_90phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1130_ _0518_ VGND VPWR _0122_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1061_ net9 VGND VPWR _0495_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_7_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0914_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ VGND VPWR _0389_ VGND VPWR sky130_fd_sc_hd__or4_2
X_0845_ _0328_ _0335_ _0337_ net69 VGND VPWR _0030_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0776_ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VPWR _0286_ VGND VPWR sky130_fd_sc_hd__and2_1
X_1259_ Dead_Time_Generator_inst_3.count_dt\[3\] Dead_Time_Generator_inst_3.count_dt\[2\]
+ _0618_ VGND VPWR _0621_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1328_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0015_ _0101_ VGND VPWR Signal_Generator_1_270phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1113_ _0517_ VGND VPWR _0106_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1044_ net12 VGND VPWR _0478_ VGND VPWR sky130_fd_sc_hd__inv_2
X_0828_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0305_ Signal_Generator_1_270phase_inst.count\[5\] VGND VPWR _0325_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0759_ _0267_ _0272_ VGND VPWR _0273_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_10_90 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1027_ _0457_ _0458_ _0459_ _0460_ VGND VPWR _0461_ VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_16_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_Dead_Time_Generator_inst_1.clk net26 VGND VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
+ VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_36 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1292_ clknet_1_0__leaf_CLK_SR _0145_ _0066_ VGND VPWR Shift_Register_Inst.data_out\[7\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1361_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0158_ VGND VPWR Dead_Time_Generator_inst_1.count_dt\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0930_ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VPWR _0401_ VGND VPWR sky130_fd_sc_hd__o31ai_1
X_0861_ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[1\]
+ VGND VPWR _0350_ VGND VPWR sky130_fd_sc_hd__and2_1
X_0792_ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR _0298_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_23_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1344_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0052_ _0117_ VGND VPWR Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1275_ _0631_ VGND VPWR _0178_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1060_ _0484_ _0491_ _0492_ _0493_ VGND VPWR _0494_ VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_0_34_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0775_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0283_ _0284_ VGND VPWR _0285_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_0844_ _0331_ _0336_ VGND VPWR _0337_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0913_ Signal_Generator_2_180phase_inst.count\[4\] net68 _0372_ _0388_ VGND VPWR
+ _0040_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_1189_ _0562_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.dt\[2\]
+ _0565_ VGND VPWR _0566_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_1258_ _0513_ _0620_ VGND VPWR _0172_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1327_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0014_ _0100_ VGND VPWR Signal_Generator_1_270phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1043_ _0469_ _0475_ _0476_ VGND VPWR _0477_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_1112_ _0446_ VGND VPWR _0517_ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_28_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0758_ Signal_Generator_1_90phase_inst.count\[2\] _0265_ VGND VPWR _0272_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0827_ Signal_Generator_1_270phase_inst.direction _0322_ _0323_ _0307_ _0324_ VGND
+ VPWR _0018_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_0689_ Shift_Register_Inst.shift_state\[2\] _0200_ Shift_Register_Inst.shift_state\[3\]
+ VGND VPWR _0221_ VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_19_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1026_ Dead_Time_Generator_inst_1.dt\[4\] Dead_Time_Generator_inst_4.count_dt\[4\]
+ VGND VPWR _0460_ VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_0_39_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1009_ _0449_ VGND VPWR _0071_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1360_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0047_ _0133_ VGND VPWR Signal_Generator_2_270phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1291_ clknet_1_0__leaf_CLK_SR _0144_ _0065_ VGND VPWR Shift_Register_Inst.data_out\[8\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0860_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0347_ _0348_ VGND VPWR _0349_ VGND VPWR sky130_fd_sc_hd__o31a_2
X_0791_ _0287_ VGND VPWR _0297_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1343_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0051_ _0116_ VGND VPWR Signal_Generator_2_90phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
X_1274_ _0513_ _0629_ _0630_ VGND VPWR _0631_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0989_ _0429_ _0436_ _0440_ _0445_ VGND VPWR net25 VGND VPWR sky130_fd_sc_hd__a31o_4
X_0912_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0368_ Signal_Generator_2_180phase_inst.count\[5\] VGND VPWR _0388_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0843_ Signal_Generator_2_0phase_inst.count\[2\] _0329_ VGND VPWR _0336_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0774_ Signal_Generator_1_180phase_inst.direction VGND VPWR _0284_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1326_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0020_ _0099_ VGND VPWR Signal_Generator_1_270phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1188_ Dead_Time_Generator_inst_1.count_dt\[2\] VGND VPWR _0565_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1257_ net62 _0618_ VGND VPWR _0620_ VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1111_ _0516_ VGND VPWR _0105_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1042_ _0470_ _0474_ VGND VPWR _0476_ VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_45_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_0757_ Signal_Generator_1_90phase_inst.count\[2\] _0268_ VGND VPWR _0271_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0826_ Signal_Generator_1_270phase_inst.count\[4\] _0305_ VGND VPWR _0324_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0688_ _0220_ VGND VPWR _0143_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1309_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0003_ _0082_ VGND VPWR Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_102 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1025_ Dead_Time_Generator_inst_4.count_dt\[4\] Dead_Time_Generator_inst_1.dt\[4\]
+ VGND VPWR _0459_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0809_ net35 VGND VPWR _0014_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_31_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_68 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0449_ VGND VPWR _0070_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1290_ clknet_1_1__leaf_CLK_SR _0143_ _0064_ VGND VPWR Shift_Register_Inst.data_out\[9\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_0790_ _0283_ _0295_ VGND VPWR _0296_ VGND VPWR sky130_fd_sc_hd__nand2_1
X_1273_ Dead_Time_Generator_inst_4.count_dt\[2\] _0626_ VGND VPWR _0630_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
X_1342_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0050_ _0115_ VGND VPWR Signal_Generator_2_90phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_0988_ _0431_ Shift_Register_Inst.data_out\[10\] _0442_ _0444_ VGND VPWR _0445_ VGND
+ VPWR sky130_fd_sc_hd__a31o_4
X_0842_ Signal_Generator_2_0phase_inst.count\[2\] _0332_ VGND VPWR _0335_ VGND VPWR
+ sky130_fd_sc_hd__xor2_1
X_0911_ net51 _0385_ _0386_ _0370_ _0387_ VGND VPWR _0039_ VGND VPWR sky130_fd_sc_hd__a32o_1
X_0773_ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ Signal_Generator_1_180phase_inst.count\[1\] Signal_Generator_1_180phase_inst.count\[0\]
+ VGND VPWR _0283_ VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_0_11_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1256_ _0513_ _0618_ _0619_ VGND VPWR _0171_ VGND VPWR sky130_fd_sc_hd__nor3_1
X_1325_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0012_ _0098_ VGND VPWR Signal_Generator_1_180phase_inst.count\[5\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1187_ _0562_ Dead_Time_Generator_inst_1.dt\[1\] _0563_ Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VPWR _0564_ VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_0_6_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1110_ _0516_ VGND VPWR _0104_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_29_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1041_ _0470_ _0474_ _0468_ _0462_ VGND VPWR _0475_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0825_ Signal_Generator_1_270phase_inst.count\[4\] _0309_ VGND VPWR _0323_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_9_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0687_ _0182_ Shift_Register_Inst.data_out\[9\] _0219_ VGND VPWR _0220_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
X_0756_ _0027_ _0269_ _0270_ VGND VPWR _0022_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1239_ Dead_Time_Generator_inst_3.count_dt\[1\] VGND VPWR _0604_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1308_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0002_ _0081_ VGND VPWR Signal_Generator_1_0phase_inst.count\[2\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_114 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1024_ Dead_Time_Generator_inst_4.count_dt\[3\] Dead_Time_Generator_inst_1.dt\[3\]
+ VGND VPWR _0458_ VGND VPWR sky130_fd_sc_hd__and2b_1
X_0808_ _0307_ _0310_ VGND VPWR _0020_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_0739_ Signal_Generator_1_0phase_inst.count\[4\] _0244_ VGND VPWR _0258_ VGND VPWR
+ sky130_fd_sc_hd__or2_1
XFILLER_0_39_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_106 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_128 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1007_ _0449_ VGND VPWR _0069_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_CLK_SR clknet_0_CLK_SR VGND VPWR clknet_1_0__leaf_CLK_SR VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1272_ Dead_Time_Generator_inst_4.count_dt\[2\] _0626_ VGND VPWR _0629_ VGND VPWR
+ sky130_fd_sc_hd__nand2_1
X_1341_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0049_ _0114_ VGND VPWR Signal_Generator_2_90phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0987_ _0439_ Shift_Register_Inst.data_out\[12\] _0443_ VGND VPWR _0444_ VGND VPWR
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0910_ Signal_Generator_2_180phase_inst.count\[4\] _0368_ VGND VPWR _0387_ VGND VPWR
+ sky130_fd_sc_hd__xnor2_1
X_0841_ _0034_ _0333_ _0334_ VGND VPWR _0029_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_0772_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0266_ _0282_ VGND VPWR _0026_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_1186_ Dead_Time_Generator_inst_1.count_dt\[0\] VGND VPWR _0563_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1255_ net50 _0616_ VGND VPWR _0619_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1324_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0011_ _0097_ VGND VPWR Signal_Generator_1_180phase_inst.count\[4\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_0_40_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1040_ Signal_Generator_2_0phase_inst.count\[5\] _0467_ _0472_ _0473_ VGND VPWR _0474_
+ VGND VPWR sky130_fd_sc_hd__o22a_1
X_0824_ _0319_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ VGND VPWR _0322_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0755_ _0263_ _0269_ net54 VGND VPWR _0270_ VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_0686_ _0187_ _0196_ Shift_Register_Inst.shift_state\[3\] VGND VPWR _0219_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_1169_ Shift_Register_Inst.data_out\[6\] Signal_Generator_1_90phase_inst.count\[3\]
+ Shift_Register_Inst.data_out\[5\] VGND VPWR _0546_ VGND VPWR sky130_fd_sc_hd__and3b_1
X_1238_ _0561_ _0573_ VGND VPWR _0169_ VGND VPWR sky130_fd_sc_hd__nor2_1
X_1307_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0001_ _0080_ VGND VPWR Signal_Generator_1_0phase_inst.count\[1\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_1023_ _0451_ Dead_Time_Generator_inst_1.dt\[2\] _0454_ _0455_ _0456_ VGND VPWR _0457_
+ VGND VPWR sky130_fd_sc_hd__o221a_1
X_0738_ _0254_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ VGND VPWR _0257_ VGND VPWR sky130_fd_sc_hd__or3b_1
X_0807_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0309_ VGND VPWR _0310_ VGND VPWR sky130_fd_sc_hd__and3_1
X_0669_ _0182_ Dead_Time_Generator_inst_1.dt\[4\] _0206_ VGND VPWR _0207_ VGND VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1006_ _0449_ VGND VPWR _0068_ VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_246 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1340_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0055_ _0113_ VGND VPWR Signal_Generator_2_90phase_inst.direction
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_1271_ _0628_ VGND VPWR _0177_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0986_ net24 _0430_ _0432_ net19 VGND VPWR _0443_ VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_1_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0771_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0261_ Signal_Generator_1_90phase_inst.count\[5\] VGND VPWR _0282_ VGND VPWR sky130_fd_sc_hd__o31a_1
X_0840_ _0328_ _0333_ net59 VGND VPWR _0334_ VGND VPWR sky130_fd_sc_hd__a21oi_1
X_1323_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0010_ _0096_ VGND VPWR Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VPWR sky130_fd_sc_hd__dfstp_1
X_1185_ Dead_Time_Generator_inst_1.count_dt\[1\] VGND VPWR _0562_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1254_ Dead_Time_Generator_inst_3.count_dt\[1\] Dead_Time_Generator_inst_3.count_dt\[0\]
+ _0615_ VGND VPWR _0618_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_46_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0969_ _0427_ VGND VPWR net17 VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_45_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0823_ _0307_ _0318_ _0321_ net61 VGND VPWR _0017_ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0754_ _0268_ _0265_ VGND VPWR _0269_ VGND VPWR sky130_fd_sc_hd__or2_1
X_0685_ _0218_ VGND VPWR _0144_ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1306_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0000_ _0079_ VGND VPWR Signal_Generator_1_0phase_inst.count\[0\]
+ VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1099_ _0515_ VGND VPWR _0094_ VGND VPWR sky130_fd_sc_hd__inv_2
X_1168_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VPWR _0545_ VGND VPWR sky130_fd_sc_hd__and3_1
X_1237_ net31 _0601_ _0561_ VGND VPWR _0168_ VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_42_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1022_ Dead_Time_Generator_inst_1.dt\[3\] Dead_Time_Generator_inst_4.count_dt\[3\]
+ VGND VPWR _0456_ VGND VPWR sky130_fd_sc_hd__or2b_1
X_0668_ _0205_ _0186_ Shift_Register_Inst.shift_state\[2\] VGND VPWR _0206_ VGND VPWR
+ sky130_fd_sc_hd__or3b_1
X_0737_ _0242_ _0253_ _0256_ Signal_Generator_1_0phase_inst.direction VGND VPWR _0003_
+ VGND VPWR sky130_fd_sc_hd__a22o_1
X_0806_ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ _0308_ VGND VPWR _0309_ VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_0_21_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold40 Signal_Generator_2_0phase_inst.count\[4\] VGND VPWR net65 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_1005_ _0449_ VGND VPWR _0067_ VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_44_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
.ends

.subckt nmos_waffle_14x14 dw_n6950_n7050# a_n938_0# a_13362_0# a_n1100_n1200#
Xnmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_0 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_1 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_source_frame_lt_10 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_rb_2 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_source_frame_lt_11 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_3 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_4 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_5 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_0 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_6 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_1 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_7 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_2 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_8 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_in_0 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_3 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_9 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_in_1 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_70 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_4 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_in_2 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_60 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_71 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_5 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_in_3 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_50 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_61 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_6 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_in_4 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_40 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_51 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_62 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_7 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_5 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_30 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_41 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_52 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_63 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_8 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_6 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_20 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_31 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_42 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_53 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_64 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_9 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_7 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_10 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_21 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_32 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_43 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_54 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_65 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_8 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_11 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_22 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_33 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_44 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_55 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_66 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_9 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_12 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_23 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_34 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_45 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_56 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_67 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_frame_lt_10 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_11 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_13362_0#
+ a_n1100_n1200# a_n938_0# a_13362_0# a_13362_0# nmos_drain_frame_lt
Xnmos_drain_in_13 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_24 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_35 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_46 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_57 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_68 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_0 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_rb_10 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_in_14 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_25 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_36 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_47 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_58 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_69 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_1 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_11 a_13362_0# a_13362_0# a_13362_0# a_13362_0# a_n938_0# a_13362_0#
+ a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# a_13362_0# nmos_drain_frame_rb
Xnmos_drain_in_15 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_26 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_37 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_48 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_59 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_2 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_16 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_27 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_38 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_49 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_3 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_17 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_28 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_39 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_4 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_18 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_drain_in_29 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_5 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_19 a_13362_0# a_13362_0# a_13362_0# dw_n6950_n7050# a_13362_0# a_13362_0#
+ a_n938_0# a_13362_0# a_13362_0# a_n1100_n1200# a_13362_0# a_13362_0# nmos_drain_in
Xnmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_6 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_7 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_8 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_9 a_n938_0# a_n938_0# a_n938_0# a_13362_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_13362_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
X0 a_13362_0# a_n1100_n1200# a_n938_0# a_13362_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X1 a_n938_0# a_n1100_n1200# a_13362_0# a_13362_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_13362_0# a_n1100_n1200# a_n938_0# a_13362_0# sky130_fd_pr__nfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_13362_0# a_13362_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt pmos_waffle_26x26 a_n1100_n1200# a_26562_0# a_n938_0#
Xpmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_230 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_frame_lt_18 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_285 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_274 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_263 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_252 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_241 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_20 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_31 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_42 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_53 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_64 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_75 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_86 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_97 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_220 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_231 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_286 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_275 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_264 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_253 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_242 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_frame_lt_19 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_10 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_21 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_32 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_43 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_54 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_65 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_76 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_87 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_98 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_210 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_221 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_232 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_254 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_243 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_287 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_276 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_265 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_11 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_22 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_33 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_44 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_55 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_66 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_77 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_88 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_99 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_in_200 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_211 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_222 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_233 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_277 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_266 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_255 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_244 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_12 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_23 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_34 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_45 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_56 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_67 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_78 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_89 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_201 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_212 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_223 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_234 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_278 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_267 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_256 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_245 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_13 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_24 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_35 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_46 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_57 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_68 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_79 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_202 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_213 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_224 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_235 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_279 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_268 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_257 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_246 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_14 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_25 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_36 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_47 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_58 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_69 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_203 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_214 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_225 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_236 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_269 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_258 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_247 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_15 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_26 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_37 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_48 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_59 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_204 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_215 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_226 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_237 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_259 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_248 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_16 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_27 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_38 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_49 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_205 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_216 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_227 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_238 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_249 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_17 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_28 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_39 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_206 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_217 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_228 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_239 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_18 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_29 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_207 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_218 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_229 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_19 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_208 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_219 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_209 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_190 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_180 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_191 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_170 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_181 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_192 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_160 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_171 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_182 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_193 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_0 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_150 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_161 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_172 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_183 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_194 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_rb_1 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_140 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_151 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_162 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_173 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_184 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_195 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_rb_2 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_130 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_141 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_152 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_163 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_174 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_185 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_196 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_rb_3 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_120 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_131 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_142 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_153 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_164 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_175 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_186 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_197 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_rb_4 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_110 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_121 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_132 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_143 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_154 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_165 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_176 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_187 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_198 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_20 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_rb_5 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_0 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_100 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_111 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_122 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_133 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_144 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_155 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_166 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_177 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_188 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_199 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_10 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_21 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_rb_20 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_6 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_101 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_112 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_123 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_134 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_145 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_0 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_1 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_156 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_167 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_178 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_189 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_11 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_22 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_0 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_frame_rb_10 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_21 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_7 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_1 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_2 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_102 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_113 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_124 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_135 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_146 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_157 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_168 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_179 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_12 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_frame_lt_23 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_1 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_frame_rb_11 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_22 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_2 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_frame_rb_8 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_3 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_103 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_114 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_125 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_136 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_147 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_158 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_169 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_13 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_2 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_frame_rb_12 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_rb_23 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_3 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_frame_rb_9 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_4 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_104 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_115 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_126 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_137 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_148 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_159 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_14 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_3 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_20 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_frame_rb_13 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_4 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_5 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_105 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_116 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_127 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_138 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_149 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_frame_lt_15 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_lt_4 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_21 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_10 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_frame_rb_14 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_in_106 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_117 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_128 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_139 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_5 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_6 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_16 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_5 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_22 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_11 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_90 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_rb_15 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_6 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_7 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_107 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_118 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_129 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_17 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_6 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_23 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_12 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_80 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_91 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_rb_16 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_7 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_8 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_108 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_119 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_lt_18 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_7 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_13 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_280 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_70 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_81 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_92 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_rb_17 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_8 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_drain_in_9 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_109 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_drain_frame_lt_19 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_frame_lt_8 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_281 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_270 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_frame_lt_14 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_60 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_71 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_82 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_93 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_rb_18 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_drain_frame_lt_9 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0#
+ a_n1100_n1200# a_n938_0# a_26562_0# a_26562_0# pmos_drain_frame_lt
Xpmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_9 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_source_frame_lt_15 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_282 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_271 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_260 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_50 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_61 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_72 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_83 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_94 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_frame_rb_19 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_frame_rb
Xpmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_16 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_283 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_272 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_261 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_250 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_40 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_51 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_62 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_73 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_84 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_95 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_rb
Xpmos_source_frame_lt_17 a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_frame_lt
Xpmos_drain_in_284 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_273 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_262 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_251 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_240 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_26562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# pmos_source_in
Xpmos_drain_in_30 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_41 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_52 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_63 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_74 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_85 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
Xpmos_drain_in_96 a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_26562_0# a_n938_0#
+ a_26562_0# a_26562_0# a_n1100_n1200# a_26562_0# a_26562_0# pmos_drain_in
X0 a_26562_0# a_n1100_n1200# a_n938_0# a_26562_0# sky130_fd_pr__pfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X1 a_n938_0# a_n1100_n1200# a_26562_0# a_26562_0# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_26562_0# a_n1100_n1200# a_n938_0# a_26562_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_26562_0# a_26562_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt power_stage_2 out nmos_waffle_14x14_1/dw_n6950_n7050# nmos_waffle_14x14_0/dw_n6950_n7050#
+ s4 s3 s2 s1 fc2 VP VN VSUBS fc1
Xnmos_waffle_14x14_0 nmos_waffle_14x14_0/dw_n6950_n7050# fc2 VN s4 nmos_waffle_14x14
Xnmos_waffle_14x14_1 nmos_waffle_14x14_1/dw_n6950_n7050# out fc2 s3 nmos_waffle_14x14
Xpmos_waffle_26x26_0 s2 fc1 out pmos_waffle_26x26
Xpmos_waffle_26x26_1 s1 VP fc1 pmos_waffle_26x26
.ends

.subckt converter_2 m1_2000_59000# power_stage_2_0/out power_stage_2_0/VP D4 D2 D3
+ VLS power_stage_2_0/nmos_waffle_14x14_1/dw_n6950_n7050# power_stage_2_0/fc1 power_stage_2_0/VN
+ VDD power_stage_2_0/nmos_waffle_14x14_0/dw_n6950_n7050# power_stage_2_0/fc2 D1 VSUBS
Xpower_stage_2_0 power_stage_2_0/out power_stage_2_0/nmos_waffle_14x14_1/dw_n6950_n7050#
+ power_stage_2_0/nmos_waffle_14x14_0/dw_n6950_n7050# power_stage_2_0/s4 power_stage_2_0/s3
+ power_stage_2_0/s2 power_stage_2_0/s1 power_stage_2_0/fc2 power_stage_2_0/VP power_stage_2_0/VN
+ VSUBS power_stage_2_0/fc1 power_stage_2
Xlevel_shifter_0 VDD VLS VSUBS D1 power_stage_2_0/s1 level_shifter
Xlevel_shifter_1 VDD VLS VSUBS D2 power_stage_2_0/s2 level_shifter
Xlevel_shifter_2 VDD VLS VSUBS D3 power_stage_2_0/s3 level_shifter
Xlevel_shifter_3 VDD VLS VSUBS D4 power_stage_2_0/s4 level_shifter
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xconverter_3_0 vccd2 io_in[11] io_analog[9] io_analog[3] io_analog[7] modulator_0/NMOS_PS3
+ w_323467_394837# io_analog[5] converter_3
Xconverter_1_0 io_analog[3] io_analog[3] converter_1_0/D4 converter_1_0/D2 converter_1_0/D3
+ io_analog[9] io_analog[7] io_analog[4] io_analog[3] io_analog[7] vccd2 converter_1_0/D1
+ io_analog[7] io_analog[6] io_analog[5] converter_1
Xmodulator_0 io_in[26] user_clock2 io_in[25] io_in[8] converter_1_0/D3 converter_2_0/D3
+ converter_1_0/D4 converter_2_0/D4 modulator_0/NMOS_PS3 converter_1_0/D1 converter_2_0/D1
+ converter_1_0/D2 converter_2_0/D2 modulator_0/PMOS_PS3 io_in[24] io_out[7] io_in[18]
+ io_in[19] io_in[20] io_in[21] io_in[22] io_in[23] io_in[9] io_in[10] io_in[14] io_in[15]
+ io_in[17] io_in[16] vccd2 io_analog[7] modulator
Xconverter_2_0 io_analog[7] io_analog[5] io_analog[3] converter_2_0/D4 converter_2_0/D2
+ converter_2_0/D3 io_analog[9] io_analog[3] io_analog[4] io_analog[7] vccd2 io_analog[3]
+ io_analog[6] converter_2_0/D1 io_analog[7] converter_2
R0 vssd2 io_oeb[6] sky130_fd_pr__res_generic_m3 w=2 l=1
R1 io_oeb[22] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R2 io_oeb[18] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R3 io_oeb[21] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R4 vccd2 io_oeb[3] sky130_fd_pr__res_generic_m3 w=2 l=1
R5 vccd2 io_oeb[10] sky130_fd_pr__res_generic_m3 w=2 l=1
R6 vccd2 io_oeb[8] sky130_fd_pr__res_generic_m3 w=2 l=1
R7 io_analog[3] io_analog[2] sky130_fd_pr__res_generic_m3 w=8.5 l=3.05
R8 io_oeb[16] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R9 io_oeb[17] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R10 vccd2 io_oeb[1] sky130_fd_pr__res_generic_m3 w=2 l=1
R11 vccd2 io_oeb[12] sky130_fd_pr__res_generic_m3 w=2 l=1
R12 io_oeb[25] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R13 io_oeb[15] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R14 vccd2 io_oeb[2] sky130_fd_pr__res_generic_m3 w=2 l=1
R15 vccd2 io_oeb[13] sky130_fd_pr__res_generic_m3 w=2 l=1
R16 vccd2 io_oeb[11] sky130_fd_pr__res_generic_m3 w=2 l=1
R17 io_oeb[20] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R18 io_oeb[24] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R19 io_oeb[19] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R20 vssd2 io_oeb[7] sky130_fd_pr__res_generic_m3 w=2 l=1
R21 io_analog[8] io_analog[7] sky130_fd_pr__res_generic_m3 w=12.5 l=3.46
R22 io_oeb[14] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R23 vccd2 io_oeb[9] sky130_fd_pr__res_generic_m3 w=2 l=1
R24 io_oeb[26] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R25 vccd2 io_oeb[4] sky130_fd_pr__res_generic_m3 w=2 l=1
R26 vccd2 io_oeb[0] sky130_fd_pr__res_generic_m3 w=2 l=1
R27 io_oeb[23] vccd2 sky130_fd_pr__res_generic_m3 w=2 l=1
R28 vccd2 io_oeb[5] sky130_fd_pr__res_generic_m3 w=2 l=1
.ends

